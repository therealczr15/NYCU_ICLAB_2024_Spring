//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2024 Spring
//   Lab01 Exercise   : Code Calculator
//   Author           : Jhan-Yi LIAO
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : CC.v
//   Module Name : CC
//   Release version : V1.0 (Release Date: 2024-02)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module CC(
  // Input signals
    opt,
    in_n0, in_n1, in_n2, in_n3, in_n4,  
  // Output signals
    out_n
);

//================================================================
//   INPUT AND OUTPUT DECLARATION                         
//================================================================
input [3:0] in_n0, in_n1, in_n2, in_n3, in_n4;
input [2:0] opt;
output reg [9:0] out_n;                  

//================================================================
//    Wire & Registers 
//================================================================
// Declare the wire/reg you would use in your circuit
// remember 
// wire for port connection and cont. assignment
// reg for proc. assignment
reg [3:0] sort[0:17];
reg [4:0] avg1;
reg signed [4:0] norm[0:4], mul1, mul2;
reg signed [8:0] mul;
reg signed [7:0] add1;
reg signed [9:0] eq1;
reg signed [9:0] add2;
reg signed [4:0] avg2;
reg signed [9:0] eq2;

//================================================================
//    DESIGN
//================================================================

CMP c1(.a(in_n0),    .b(in_n3),    .s(sort[0]),  .l(sort[1]));
CMP c2(.a(in_n1),    .b(in_n4),    .s(sort[2]),  .l(sort[3]));
CMP c3(.a(sort[0]),  .b(in_n2),    .s(sort[4]),  .l(sort[5]));
CMP c4(.a(sort[2]),  .b(sort[1]),  .s(sort[6]),  .l(sort[7]));
CMP c5(.a(sort[4]),  .b(sort[6]),  .s(sort[8]),  .l(sort[9]));
CMP c6(.a(sort[5]),  .b(sort[3]),  .s(sort[10]), .l(sort[11]));
CMP c7(.a(sort[9]),  .b(sort[10]), .s(sort[12]), .l(sort[13]));
CMP c8(.a(sort[7]),  .b(sort[11]), .s(sort[14]), .l(sort[15]));
CMP c9(.a(sort[13]), .b(sort[14]), .s(sort[16]), .l(sort[17]));

always @(*) begin
  if(opt[0]) begin
    avg1 = (sort[8] + sort[15]) >> 1;
  end
  else begin
    avg1 = 0;
  end
end

always @(*) begin
  if(!opt[1]) begin
    norm[0] = sort[8]  - avg1;
    norm[1] = sort[12] - avg1;
    norm[2] = sort[16] - avg1;
    norm[3] = sort[17] - avg1;
    norm[4] = sort[15] - avg1;
  end
  else begin
    norm[0] = sort[15] - avg1;
    norm[1] = sort[17] - avg1;
    norm[2] = sort[16] - avg1;
    norm[3] = sort[12] - avg1;
    norm[4] = sort[8]  - avg1;
  end
end

always @(*) begin
  if(opt[2]) begin
    mul1 = norm[0];
    mul2 = norm[4];
  end
  else begin
    mul1 = norm[1];
    mul2 = norm[2];
  end
end

always @(*) begin
  mul = mul1 * mul2;
  add1 = ((norm[0] + norm[1]) + norm[2] + (norm[3] + norm[4]));
  eq1 = norm[3] * 3 - mul;
  add2 = ((norm[0] + mul) + avg2 * norm[3]);
end

always @(*) begin
  case(add1)
    -8'd19:  avg2 = -3;  -8'd18:  avg2 = -3;  -8'd17: avg2 = -3;  -8'd16: avg2 = -3;
    -8'd15:  avg2 = -3;  -8'd14:  avg2 = -2;  -8'd13: avg2 = -2;  -8'd12: avg2 = -2; -8'd11:  avg2 = -2;
    -8'd10:  avg2 = -2;  -8'd9:   avg2 = -1;  -8'd8:  avg2 = -1;  -8'd7:  avg2 = -1; -8'd6:   avg2 = -1;
    -8'd5:   avg2 = -1;  -8'd4:   avg2 =  0;  -8'd3:  avg2 =  0;  -8'd2:  avg2 =  0; -8'd1:   avg2 =  0; 
     8'd0:   avg2 =  0;   8'd1:   avg2 =  0;   8'd2:  avg2 =  0;   8'd3:  avg2 =  0;  8'd4:   avg2 =  0;
     8'd5:   avg2 =  1;   8'd6:   avg2 =  1;   8'd7:  avg2 =  1;   8'd8:  avg2 =  1;  8'd9:   avg2 =  1;
     8'd10:  avg2 =  2;   8'd11:  avg2 =  2;   8'd12: avg2 =  2;   8'd13: avg2 =  2;  8'd14:  avg2 =  2;
     8'd15:  avg2 =  3;   8'd16:  avg2 =  3;   8'd17: avg2 =  3;   8'd18: avg2 =  3;  8'd19:  avg2 =  3;
     8'd20:  avg2 =  4;   8'd21:  avg2 =  4;   8'd22: avg2 =  4;   8'd23: avg2 =  4;  8'd24:  avg2 =  4;
     8'd25:  avg2 =  5;   8'd26:  avg2 =  5;   8'd27: avg2 =  5;   8'd28: avg2 =  5;  8'd29:  avg2 =  5;
     8'd30:  avg2 =  6;   8'd31:  avg2 =  6;   8'd32: avg2 =  6;   8'd33: avg2 =  6;  8'd34:  avg2 =  6;
     8'd35:  avg2 =  7;   8'd36:  avg2 =  7;   8'd37: avg2 =  7;   8'd38: avg2 =  7;  8'd39:  avg2 =  7;
     8'd40:  avg2 =  8;   8'd41:  avg2 =  8;   8'd42: avg2 =  8;   8'd43: avg2 =  8;  8'd44:  avg2 =  8;
     8'd45:  avg2 =  9;   8'd46:  avg2 =  9;   8'd47: avg2 =  9;   8'd48: avg2 =  9;  8'd49:  avg2 =  9;
     8'd50:  avg2 =  10;  8'd51:  avg2 =  10;  8'd52: avg2 =  10;  8'd53: avg2 =  10; 8'd54:  avg2 =  10;
     8'd55:  avg2 =  11;  8'd56:  avg2 =  11;  8'd57: avg2 =  11;  8'd58: avg2 =  11; 8'd59:  avg2 =  11;
     8'd60:  avg2 =  12;  8'd61:  avg2 =  12;  8'd62: avg2 =  12;  8'd63: avg2 =  12; 8'd64:  avg2 =  12;
     8'd65:  avg2 =  13;  8'd66:  avg2 =  13;  8'd67: avg2 =  13;  8'd68: avg2 =  13; default : avg2 = 0;
  endcase
end

always @(*) begin
  case(add2)
    -10'd50:  eq2 = -16; -10'd49:  eq2 = -16; -10'd48:  eq2 = -16;
    -10'd47:  eq2 = -15; -10'd46:  eq2 = -15; -10'd45:  eq2 = -15;
    -10'd44:  eq2 = -14; -10'd43:  eq2 = -14; -10'd42:  eq2 = -14;
    -10'd41:  eq2 = -13; -10'd40:  eq2 = -13; -10'd39:  eq2 = -13;
    -10'd38:  eq2 = -12; -10'd37:  eq2 = -12; -10'd36:  eq2 = -12;
    -10'd35:  eq2 = -11; -10'd34:  eq2 = -11; -10'd33:  eq2 = -11;
    -10'd32:  eq2 = -10; -10'd31:  eq2 = -10; -10'd30:  eq2 = -10;
    -10'd29:  eq2 = -9;  -10'd28:  eq2 = -9;  -10'd27:  eq2 = -9;
    -10'd26:  eq2 = -8;  -10'd25:  eq2 = -8;  -10'd24:  eq2 = -8;
    -10'd23:  eq2 = -7;  -10'd22:  eq2 = -7;  -10'd21:  eq2 = -7;
    -10'd20:  eq2 = -6;  -10'd19:  eq2 = -6;  -10'd18:  eq2 = -6;
    -10'd17:  eq2 = -5;  -10'd16:  eq2 = -5;  -10'd15:  eq2 = -5;
    -10'd14:  eq2 = -4;  -10'd13:  eq2 = -4;  -10'd12:  eq2 = -4;
    -10'd11:  eq2 = -3;  -10'd10:  eq2 = -3;  -10'd9:   eq2 = -3;
    -10'd8:   eq2 = -2;  -10'd7:   eq2 = -2;  -10'd6:   eq2 = -2;
    -10'd5:   eq2 = -1;  -10'd4:   eq2 = -1;  -10'd3:   eq2 = -1;
    -10'd2:   eq2 =  0;  -10'd1:   eq2 =  0;   10'd0:   eq2 =  0;
     10'd1:   eq2 =  0;   10'd2:   eq2 =  0;   
     10'd3:   eq2 =  1;   10'd4:   eq2 =  1;   10'd5:   eq2 =  1;   
     10'd6:   eq2 =  2;   10'd7:   eq2 =  2;   10'd8:   eq2 =  2;
     10'd9:   eq2 =  3;   10'd10:  eq2 =  3;   10'd11:  eq2 =  3;
     10'd12:  eq2 =  4;   10'd13:  eq2 =  4;   10'd14:  eq2 =  4;
     10'd15:  eq2 =  5;   10'd16:  eq2 =  5;   10'd17:  eq2 =  5;
     10'd18:  eq2 =  6;   10'd19:  eq2 =  6;   10'd20:  eq2 =  6;
     10'd21:  eq2 =  7;   10'd22:  eq2 =  7;   10'd23:  eq2 =  7;
     10'd24:  eq2 =  8;   10'd25:  eq2 =  8;   10'd26:  eq2 =  8;
     10'd27:  eq2 =  9;   10'd28:  eq2 =  9;   10'd29:  eq2 =  9;
     10'd30:  eq2 =  10;  10'd31:  eq2 =  10;  10'd32:  eq2 =  10;
     10'd33:  eq2 =  11;  10'd34:  eq2 =  11;  10'd35:  eq2 =  11;
     10'd36:  eq2 =  12;  10'd37:  eq2 =  12;  10'd38:  eq2 =  12;
     10'd39:  eq2 =  13;  10'd40:  eq2 =  13;  10'd41:  eq2 =  13;
     10'd42:  eq2 =  14;  10'd43:  eq2 =  14;  10'd44:  eq2 =  14;
     10'd45:  eq2 =  15;  10'd46:  eq2 =  15;  10'd47:  eq2 =  15;
     10'd48:  eq2 =  16;  10'd49:  eq2 =  16;  10'd50:  eq2 =  16;
     10'd51:  eq2 =  17;  10'd52:  eq2 =  17;  10'd53:  eq2 =  17;
     10'd54:  eq2 =  18;  10'd55:  eq2 =  18;  10'd56:  eq2 =  18;
     10'd57:  eq2 =  19;  10'd58:  eq2 =  19;  10'd59:  eq2 =  19;
     10'd60:  eq2 =  20;  10'd61:  eq2 =  20;  10'd62:  eq2 =  20;
     10'd63:  eq2 =  21;  10'd64:  eq2 =  21;  10'd65:  eq2 =  21;
     10'd66:  eq2 =  22;  10'd67:  eq2 =  22;  10'd68:  eq2 =  22;
     10'd69:  eq2 =  23;  10'd70:  eq2 =  23;  10'd71:  eq2 =  23;
     10'd72:  eq2 =  24;  10'd73:  eq2 =  24;  10'd74:  eq2 =  24;
     10'd75:  eq2 =  25;  10'd76:  eq2 =  25;  10'd77:  eq2 =  25;
     10'd78:  eq2 =  26;  10'd79:  eq2 =  26;  10'd80:  eq2 =  26;
     10'd81:  eq2 =  27;  10'd82:  eq2 =  27;  10'd83:  eq2 =  27;
     10'd84:  eq2 =  28;  10'd85:  eq2 =  28;  10'd86:  eq2 =  28;
     10'd87:  eq2 =  29;  10'd88:  eq2 =  29;  10'd89:  eq2 =  29;
     10'd90:  eq2 =  30;  10'd91:  eq2 =  30;  10'd92:  eq2 =  30;
     10'd93:  eq2 =  31;  10'd94:  eq2 =  31;  10'd95:  eq2 =  31;
     10'd96:  eq2 =  32;  10'd97:  eq2 =  32;  10'd98:  eq2 =  32;
     10'd99:  eq2 =  33;  10'd100: eq2 =  33;  10'd101: eq2 =  33;
     10'd102: eq2 =  34;  10'd103: eq2 =  34;  10'd104: eq2 =  34;
     10'd105: eq2 =  35;  10'd106: eq2 =  35;  10'd107: eq2 =  35;
     10'd108: eq2 =  36;  10'd109: eq2 =  36;  10'd110: eq2 =  36;
     10'd111: eq2 =  37;  10'd112: eq2 =  37;  10'd113: eq2 =  37;
     10'd114: eq2 =  38;  10'd115: eq2 =  38;  10'd116: eq2 =  38;
     10'd117: eq2 =  39;  10'd118: eq2 =  39;  10'd119: eq2 =  39;
     10'd120: eq2 =  40;  10'd121: eq2 =  40;  10'd122: eq2 =  40;
     10'd123: eq2 =  41;  10'd124: eq2 =  41;  10'd125: eq2 =  41;
     10'd126: eq2 =  42;  10'd127: eq2 =  42;  10'd128: eq2 =  42;
     10'd129: eq2 =  43;  10'd130: eq2 =  43;  10'd131: eq2 =  43;
     10'd132: eq2 =  44;  10'd133: eq2 =  44;  10'd134: eq2 =  44;
     10'd135: eq2 =  45;  10'd136: eq2 =  45;  10'd137: eq2 =  45;
     10'd138: eq2 =  46;  10'd139: eq2 =  46;  10'd140: eq2 =  46;
     10'd141: eq2 =  47;  10'd142: eq2 =  47;  10'd143: eq2 =  47;
     10'd144: eq2 =  48;  10'd145: eq2 =  48;  10'd146: eq2 =  48;
     10'd147: eq2 =  49;  10'd148: eq2 =  49;  10'd149: eq2 =  49;
     10'd150: eq2 =  50;  10'd151: eq2 =  50;  10'd152: eq2 =  50;
     10'd153: eq2 =  51;  10'd154: eq2 =  51;  10'd155: eq2 =  51;
     10'd156: eq2 =  52;  10'd157: eq2 =  52;  10'd158: eq2 =  52;
     10'd159: eq2 =  53;  10'd160: eq2 =  53;  10'd161: eq2 =  53;
     10'd162: eq2 =  54;  10'd163: eq2 =  54;  10'd164: eq2 =  54;
     10'd165: eq2 =  55;  10'd166: eq2 =  55;  10'd167: eq2 =  55;
     10'd168: eq2 =  56;  10'd169: eq2 =  56;  10'd170: eq2 =  56;
     10'd171: eq2 =  57;  10'd172: eq2 =  57;  10'd173: eq2 =  57;
     10'd174: eq2 =  58;  10'd175: eq2 =  58;  10'd176: eq2 =  58;
     10'd177: eq2 =  59;  10'd178: eq2 =  59;  10'd179: eq2 =  59;
     10'd180: eq2 =  60;  10'd181: eq2 =  60;  10'd182: eq2 =  60;
     10'd183: eq2 =  61;  10'd184: eq2 =  61;  10'd185: eq2 =  61;
     10'd186: eq2 =  62;  10'd187: eq2 =  62;  10'd188: eq2 =  62;
     10'd189: eq2 =  63;  10'd190: eq2 =  63;  10'd191: eq2 =  63;
     10'd192: eq2 =  64;  10'd193: eq2 =  64;  10'd194: eq2 =  64;
     10'd195: eq2 =  65;  10'd196: eq2 =  65;  10'd197: eq2 =  65;
     10'd198: eq2 =  66;  10'd199: eq2 =  66;  10'd200: eq2 =  66;
     10'd201: eq2 =  67;  10'd202: eq2 =  67;  10'd203: eq2 =  67;
     10'd204: eq2 =  68;  10'd205: eq2 =  68;  10'd206: eq2 =  68;
     10'd207: eq2 =  69;  10'd208: eq2 =  69;  10'd209: eq2 =  69;
     10'd210: eq2 =  70;  10'd211: eq2 =  70;  10'd212: eq2 =  70;
     10'd213: eq2 =  71;  10'd214: eq2 =  71;  10'd215: eq2 =  71;
     10'd216: eq2 =  72;  10'd217: eq2 =  72;  10'd218: eq2 =  72;
     10'd219: eq2 =  73;  10'd220: eq2 =  73;  10'd221: eq2 =  73;
     10'd222: eq2 =  74;  10'd223: eq2 =  74;  10'd224: eq2 =  74;
     10'd225: eq2 =  75;  10'd226: eq2 =  75;  10'd227: eq2 =  75;
     10'd228: eq2 =  76;  10'd229: eq2 =  76;  10'd230: eq2 =  76;
     10'd231: eq2 =  77;  10'd232: eq2 =  77;  10'd233: eq2 =  77;
     10'd234: eq2 =  78;  10'd235: eq2 =  78;  10'd236: eq2 =  78;
     10'd237: eq2 =  79;  10'd238: eq2 =  79;  10'd239: eq2 =  79;
     10'd240: eq2 =  80;  10'd241: eq2 =  80;  10'd242: eq2 =  80;
     10'd243: eq2 =  81;  10'd244: eq2 =  81;  10'd245: eq2 =  81;
     10'd246: eq2 =  82;  10'd247: eq2 =  82;  10'd248: eq2 =  82;
     10'd249: eq2 =  83;  10'd250: eq2 =  83;  10'd251: eq2 =  83;
     10'd252: eq2 =  84;  10'd253: eq2 =  84;  10'd254: eq2 =  84;
     10'd255: eq2 =  85;  10'd256: eq2 =  85;  10'd257: eq2 =  85;
     10'd258: eq2 =  86;  10'd259: eq2 =  86;  10'd260: eq2 =  86;
     10'd261: eq2 =  87;  10'd262: eq2 =  87;  10'd263: eq2 =  87;
     10'd264: eq2 =  88;  10'd265: eq2 =  88;  10'd266: eq2 =  88;
     10'd267: eq2 =  89;  10'd268: eq2 =  89;  10'd269: eq2 =  89;
     10'd270: eq2 =  90;  10'd271: eq2 =  90;  10'd272: eq2 =  90;
     10'd273: eq2 =  91;  10'd274: eq2 =  91;  10'd275: eq2 =  91;
     10'd276: eq2 =  92;  10'd277: eq2 =  92;  10'd278: eq2 =  92;
     10'd279: eq2 =  93;  10'd280: eq2 =  93;  10'd281: eq2 =  93;
     10'd282: eq2 =  94;  10'd283: eq2 =  94;  10'd284: eq2 =  94;
     10'd285: eq2 =  95;  10'd286: eq2 =  95;  10'd287: eq2 =  95;
     10'd288: eq2 =  96;  10'd289: eq2 =  96;  10'd290: eq2 =  96;
     10'd291: eq2 =  97;  10'd292: eq2 =  97;  10'd293: eq2 =  97;
     10'd294: eq2 =  98;  10'd295: eq2 =  98;  10'd296: eq2 =  98;
     10'd297: eq2 =  99;  10'd298: eq2 =  99;  10'd299: eq2 =  99;
     10'd300: eq2 =  100; 10'd301: eq2 =  100; 10'd302: eq2 =  100;
     10'd303: eq2 =  101; 10'd304: eq2 =  101; 10'd305: eq2 =  101;
     10'd306: eq2 =  102; 10'd307: eq2 =  102; 10'd308: eq2 =  102;
     10'd309: eq2 =  103; 10'd310: eq2 =  103; 10'd311: eq2 =  103;
     10'd312: eq2 =  104; 10'd313: eq2 =  104; 10'd314: eq2 =  104;
     10'd315: eq2 =  105; 10'd316: eq2 =  105; 10'd317: eq2 =  105;
     10'd318: eq2 =  106; 10'd319: eq2 =  106; 10'd320: eq2 =  106;
     10'd321: eq2 =  107; 10'd322: eq2 =  107; 10'd323: eq2 =  107;
     10'd324: eq2 =  108; 10'd325: eq2 =  108; 10'd326: eq2 =  108;
     10'd327: eq2 =  109; 10'd328: eq2 =  109; 10'd329: eq2 =  109;
     10'd330: eq2 =  110; 10'd331: eq2 =  110; 10'd332: eq2 =  110;
     10'd333: eq2 =  111; 10'd334: eq2 =  111; 10'd335: eq2 =  111;
     10'd336: eq2 =  112; 10'd337: eq2 =  112; 10'd338: eq2 =  112;
     10'd339: eq2 =  113; 10'd340: eq2 =  113; 10'd341: eq2 =  113;
     10'd342: eq2 =  114; 10'd343: eq2 =  114; 10'd344: eq2 =  114;
     10'd345: eq2 =  115; 10'd346: eq2 =  115; 10'd347: eq2 =  115;
     10'd348: eq2 =  116; 10'd349: eq2 =  116; 10'd350: eq2 =  116;
     10'd351: eq2 =  117; 10'd352: eq2 =  117; 10'd353: eq2 =  117;
     10'd354: eq2 =  118; 10'd355: eq2 =  118; 10'd356: eq2 =  118;
     10'd357: eq2 =  119; 10'd358: eq2 =  119; 10'd359: eq2 =  119;
     10'd360: eq2 =  120; 10'd361: eq2 =  120; 10'd362: eq2 =  120;
     10'd363: eq2 =  121; 10'd364: eq2 =  121; 10'd365: eq2 =  121;
     10'd366: eq2 =  122; 10'd367: eq2 =  122; 10'd368: eq2 =  122;
     10'd369: eq2 =  123; 10'd370: eq2 =  123; 10'd371: eq2 =  123;
     10'd372: eq2 =  124; 10'd373: eq2 =  124; 10'd374: eq2 =  124;
     10'd375: eq2 =  125; 10'd376: eq2 =  125; 10'd377: eq2 =  125;
     10'd378: eq2 =  126; 10'd379: eq2 =  126; 10'd380: eq2 =  126;
     10'd381: eq2 =  127; 10'd382: eq2 =  127; 10'd383: eq2 =  127;
     10'd384: eq2 =  128; 10'd385: eq2 =  128; 10'd386: eq2 =  128;
     10'd387: eq2 =  129; 10'd388: eq2 =  129; 10'd389: eq2 =  129;
     10'd390: eq2 =  130; 10'd391: eq2 =  130; 10'd392: eq2 =  130;
     10'd393: eq2 =  131; 10'd394: eq2 =  131; 10'd395: eq2 =  131;
     10'd396: eq2 =  132; 10'd397: eq2 =  132; 10'd398: eq2 =  132;
     10'd399: eq2 =  133; 10'd400: eq2 =  133; 10'd401: eq2 =  133;
     10'd402: eq2 =  134; 10'd403: eq2 =  134; 10'd404: eq2 =  134;
     10'd405: eq2 =  135; 10'd406: eq2 =  135; 10'd407: eq2 =  135;
     10'd408: eq2 =  136; 10'd409: eq2 =  136; 10'd410: eq2 =  136;
     10'd411: eq2 =  137; 10'd412: eq2 =  137; 10'd413: eq2 =  137;
     10'd414: eq2 =  138; 10'd415: eq2 =  138; 10'd416: eq2 =  138;
     10'd417: eq2 =  139; 10'd418: eq2 =  139; 10'd419: eq2 =  139;
     default: eq2 =  0;
  endcase
end

always @(*) begin
  if(opt[2]) begin
    if(eq1[9]) begin
      out_n = -eq1;
    end
    else begin
      out_n = eq1;
    end
  end
  else begin
    out_n = eq2;
  end
end

endmodule

//================================================================
//    Self Define Module
//================================================================
module CMP(
  // Input signals
    a, b,
  // Output signals
    s, l
);

input  [3:0] a, b;
output [3:0] s, l;

assign s = (a < b)? a : b;
assign l = (a < b)? b : a;

endmodule
