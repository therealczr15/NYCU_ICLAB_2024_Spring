//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2023 ICLAB Fall Course
//   Lab03      : BRIDGE
//   Author     : Tzu-Yun Huang
//	 Editor		: Ting-Yu Chang
//                
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : pseudo_DRAM.v
//   Module Name : pseudo_DRAM
//   Release version : v3.0 (Release Date: Sep-2023)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module pseudo_DRAM
`protected
ETg><J-4Je?<0P@J@e)J1]eTYWJC/[B,&:;?5e,515HH86eMRD;?))50a\202?g-
e(Z8/GcG0-\;]dN#YGO#1?5X5,Z9AcIfBRTRR]PM?a5;?O^(0GfHS)(5#_&/MHgF
KAPHb<66F]CYJ-9(f#Hg_:=5CRC(N3=fSCKUeADQc27NA)YM_BUFCBN_NK<\2NKB
9FGRG.]T,XFaHK/PKHXLQS7[]MT-G-&N\<EcQ1c/4?f]E\7THYOJQI&-+5R_3@dA
9]-F,S3g-2.W[D,;I#RVN8f>Y/M#@=K^[OdN(60NTCG,8M+c]SRKU#A>/,QXD)eY
&D^.W&;-UgX:b+S&4FPfRHTb4KYO&[Nb\f<YL+T(8G3(PcA40A#KZ=.K,]GTcA09
N&QK\SH8e=.2cC@(C?S8TFKSaEg,EL3Y1E3])D8(cY]fR1dXV[FORS6LVDf3Q48G
W_]9P(,KK+CM-E(M[YB#-Y@\H7F7_\eW04SL^R0SQ8J0<c8N.[6Z([3WG0VWca)G
OF+5U))UccHcI-7:J,0DV^g>@L1>-)?:a,2#@Z@dAA[Y=#1Mgg-OP0?\^bR+ScLf
[#L(R:NATC-,@PDQ^N34A3K-O3,aAGFFZM9C=NQ-B.DC35X8]Q\NXf-X3Z2\QHf;
K[DHVN4=&D\\-Q[/1^P4OfLgPK@:^N>#Dg7bHN+7?LPIET>\e]9O^N#BB,HY#GNM
fe?L(aA,(^<?=.DaV/L;-_/Hb2>&d@/J[e0c?f:7;.CPWb,]#LeP2-1YH,.?dIa^
Bb)=#PO+T]gC[:8I<G73<Sa3=)VGUG.THNBc1LB(>WH)QJ00-@H9>CQ0Td0_HcF3
RSKB2/+0ZF7gN7dS-fUXNS62TaTGDFeG26Z\,#+e^2AQ17U@d][V\2I#B3[=-:^e
NE)@^OVd#X-?LIHeO4Cd8(6(O(@Ec?;)&BZ7&J>LZMKJbZ0>ZgX&/:[IScAZ7P0U
NaG5^9-_>c_U+PQAM.WA20cR9G>RV;.1GQEZP0;3CSIW0\8@0P;J@G2c)d.UcJA(
&X5K[<.FD2F2\JWM1W5ZI9T\Z)bH=^1VK+XdYQ+A-GbX5H4?fQTHR7:W,E;(I>_7
(+J<Aa=M69I\aQg#(DaLgE4AIdbW5R(e:@)20HV0ZfV:PDZ?eW3E.fQH6H?)]Q6C
bXTZA(a7S8eHgd0]/#DJAI+DO^C>TB<fLCG/MYTD0\&H?Z&ANW=#SAT.U^9QL+_I
R^Y/\e9Z<:Y\/V4SYZ9aU^)(J2855,AP?-T7,IBc97X6>H@E9^@[180_>HJ0)69<
LD#CB&c3\RZ72aG,F[TJD[CV=T5LAW2g>Pa,G[U:YZ0(@IYD&U@L5E5T;Q36,Q7a
7T+TL+GO1N>ROIMSS.5Fa9\YZfB67)L?K&N)f3DgUVdV^dFZ4+4+Yd&7d/SK)b.=
LU&bV<5^5K6@FQP/;XGC<16^e4CAXEQS_a;C?2:3=W[E7d?RI@IC(Ea]<fA40^N3
DY\.>U[b;\cPa.&T[fOFA\8H[g\+QY71QH4D(\TBAW^UTbaa<YBB?S>Y;XR;;IQ6
dA>.[.&+b&ddUdLOS4^0YBa5aX8\eY;=^<<A63Qd5C5,]f#7XYY+7f8\(JJ0S_81
d41B>a;gX^G9PcT\U+Yf0F=EY@D[_Bc\&1#:^YWU?DW<+DNc[/>\(:PF_;5QA:A?
K,/GQFS]0J)=CNIWWV.:3.R(-_K56F7IHUG,:Kd1OV&>.CBDAT5#.\D]:KAbRJ:L
)J#[RZ--#8X<_]9#QgZ>g;3EcbMG]L9WSVRZ1(F;2(ASJK#?G1,&F?:d\>Y9X3=0
WCa<Ug0c/BOSS00OFNLN+-T)PCP-_#8;Z#AH/eBM9a##Y+ETc8&U1=&:&fMg):7C
75a26;ce>3N:^8+)b2<&-05.bPY:L)3K_I=W5@VEOV=\-a>,&[b[fU\dR._C94H;
Ec_FEWEQ13;#Y&VKWR^^B&HeYB>^4Z\LGWJE\9V41=B::V0NSdad_T;5/]gMH0GE
MB8NEGb71J1L?RMgN@L^17?AY=g&E#bT1DfW/,6P,;<.BI&c0;=E+&U8c:RS;4HH
G7)<05&TFB>D?PDG-N-1(Vb(ge.Y5)@]^6e:gU7Zb;CCZ3#+JT)A.I2L?W=6-;/5
WC<IN#B9?e-IPO3@OW=.1X.0CYIQd^5NF\^6eJ_DEUXXLFAMcdgfCbV3PY+\S28&
.^Y^.,SG=8a([cQRe(Ub=PJ>VJ<HGXE^=VM#JKc#e#ZSP:(a>6=1N.G3=](b9^E0
Pa\Te8\N-&]X5c#)BX_W(RdBPZ77<N>;g3^WKd#E2Q:L(07b20cGDOaKK^L2.f=U
?VQ3D5:CK)VD2T6RBK_Ga3fDZVIBVEL[@-S2LM<+Y7MFdaRIH1SG:^Z0F<NGYYME
_d^XK06=)>ZZg(+D_Z:5E3\L-/Q(HOEX5/5d:?&PJ9O)dYE,eSF3:(2UAV>GV9:5
JM>&cM^ELI[^C-YISGcE&7<6UJO]E4S#LAZF#O@PPd7<64)g,7JDXMVKeL^0OPD-
,ZJ3G<RccgQE>_T77/e#(ML8X8/RP5.RX3N@5=5g_I7U+_;Q>c]=HV3R4FQSg1L4
C,0B)OWSD((VedO(C.2#DM9&c(?L<FRQT;7I>V6T-<a8B&Z69(THBNW36?+WZA\(
MX?PS2g0M&[\G#<WdO.3Y@WcIZ(Y##7K29Gc_\6-\?S:@LbKg4XBUPD=SP]cB7&=
-N7FHSH><0Xb>VTM)_Nd,NYMbeVabC1^2SaF\c\8B)&<f>2N0X+N?cH/Z/L\1;K8
FN?77=?ZQ5V<A]9?^[a1_eG8ZB&IS;V]\c:[HH14Ba=[4HS,_A>K:+-:T@:FE&M3
=+LP^a:_OgeFEF?c;GO#<\Ra\BTRC_JBFOMRU2\YN]&D.=)ZLaLQBH93O,R.gZf<
Dgf7#Y=8?0=->)dIX]5Tf92OO/\HHK?aS/,a[f>D.LX2[Q-;RXWJ/aF#G:@#QMQV
Ib@;-2c-Vf.Q=>8abdF/WPGaU[OMO6Pc^HFXZ#1gCUCR9=f\FRU@X(L<N702FV=f
J5K5<B1,)WSad-H.JFVQY)I>]R2C:c5FRagCM7R>.#5V4G;T42bZde7A,((b;)Y?
@;XN\Bg1a#L7Jc73A[#W2U.4[9=NN2?+MRZa)NgGSbQC0(P>0>3<RA\bU>Z6N7ST
/@:_aSf6A=c?AE0<XA9?>>OHYE1<^,38d=,:J;c@,DO><;fQdg8^=&XP:CO_97SO
^ZM(GMB:5F,@AE-@B\DD9?WfH6=)]S1JN\,W[:/LR&O7cM;a/WYAMM#+;ZG5g8W.
I+X>#\/22I;J2]-FJ5I<1D<cdO\RHL<CZ9g1HNMR[16_,6fL\<O/75?LY1e-Geb)
)bU<Nb(cKNWFNS=F<I;DP1V.a@d6)2bd4&eUH81ZSN</)=02IGcJV\)]F5cF4\:A
f=@V;;>2:9ac#<Hd:b36dC0dJ&)XPC2Y+6C,=_:0+cXWTAe_0?<6c3#C7[UP&UJ3
EeODN>?-/>d.0,[YTHMH28\d77Mb,R90/8IQX9ge[Lb=0c0Td:5&gB[Y+9RW74?A
fBP0YG)T2AJd:;P)?7_=L8E6QAR3Qf+635)[gfDd&)#(-3_)\@)4+?UVD=4[VTPR
Gg^MZW-2IE.OOFCR^VQL/7#I)?W.XXP^Y_(EHg&_a\IBd@>GE^-D19a)edIMI[=]
b0PX;OK&WTFdJ].#Ad651ICG451RD&:&.d2ObK_H2WWP@,I[bO)3LUX3K&<1P32D
-#OaI#5RK)J]O\:=fFFL0UaUYPT1??@a9QRe&_0Y0/9E#Y</A9THg@Q/VaQPQ:Oe
7FOV+8L=30?6V#RIBVQbK.QBLOT)Z@IUObVIg3H<KIgY2(F3(aB5Z7+b[VVQ]@9U
.N5H\K#>/Ed?+L;>:9)W5A/R.V\Oa9fFLc\EK)M-e9<XMFJIeL?Y<M/V8bNYL(/T
b?Wbe#WPQ=8cG+b&B/-f>c.4JS,@H4fK>.DJR7J:)LK(2&=c3E08F#4H0O<EQ^,Y
ND_I@+Z)<31>Y<V><;4YWA4[.ZL;\>T?Q\4#XJTeGa>8;-K9NK4a)aD<):M1LD/K
8\G#GEg#>#,/8aR;.N[SA#<?+EPe,3TM\/3g)2(604-K47^2XKae)+BNXbaTL2Z/
f<?#e8THY@#C@dP+OBGZQU?7DKMN0W=<8TYZ-H<?+_e:-ZfL,H7RQPM7&ZHAV\>@
=A..BY4P+U2^OCfR1_B<d:<[f0^DL(RD(#P@e=-(Ga>ORg\#dV2U7ZD,R+&?L)LJ
+-AP;-M8:g5IR5([8K,Q8M3??0_GJ-HGc/a[O#UXNBVA242P&W@:L<+4c<gF:;S]
\\&SbeV_^e9,_dE0^9GO@Ld.YKS-4LOO_5Q6G/Aae[8eUEH?SQRHN1gF+JcEEWM+
KbCI9B&c)EWOdc(<&a_@6+214>+G7S@:#\HJXMYDM^4E=X,.SQfO,G)-MeHGP,9A
Q,Qe9DX[H+.VL/>]f5AG?c,QJ?&0W@VX@^EAW58G91bMbJ7DA8RS(30?H8N0\DIY
&d=]5]B:;W;f6P=(9\#0,OVCNb::C@_[W/U&^)Y@Z616fIWWY&9#\_P]BLJX6CVF
0T9PE_M\#e2C_Tg30HV>8=RC2.2D^<=[WfIPO5W@3M;;1c/:^eM\G0,FN\8&E<BE
PaJ^8:HUe^GdX]/O^0-9LMc:bTVIS7ZgcMJ-=QTH75fYF/f]Aa?@eN(Ob,;W^dD6
@3:JV;YXRNL7dc,<B&S#KaI[6Og,W2PE[Q?)DYPHbPW/<2aSA,6P)d:X09c@2A9b
DNR[MgKUJb9)T>07BN.DG@T^K(:-]P;gYMET8AJKPGRF:gTCAdQa^Z[M.b&1fEU@
Ked1)]65O_,ZHN4OFJ=#RdEFT3U<IX0[)<#P^IWdJ;1G:eHR@U/)7PZP53AXfH5#
04RD._cA=c5W.JG.3<71bd^HOSceeIC4#PXF?V_ZBT:<V5aT6NIQ@33@E&EEE0ZW
g_e&0#9@]O9+<.[;+#W>67SKWaDH?ATR>^W\?Bc</dAS<<QQ&#?Z]SD0OBKUF=N4
H=72T9VbSQP^N@068WF)G(&P+f.=60C.M2\IPDR;J)Z)eg[6+GFAH+J,dO)U\1_,
;=,D#VK12\>0Q3@8f^.RY?4.F[;G)6<gV@\XOe5>)(-+.BcY70gZeKYcA;PBRCHH
DbG]1F+&JKRLSEX\DC;;ECeKfcLL_WNXS7E5<dJJ@380J;f@LFf_1P-9W?I/ZcCK
(_Vfa7@:#fX?]XBS#TVCgYH^[2gEgW0:)(G)]Q1da5&O[/=TTS1b>+R)FG:TD?I)
5>N>-A]R^RR.+X[DJH=FI;7LUGI,>(5@/3RFCR,-M>5cYCAHcYT<JT7RQQ9ZJQJQ
QXANG5-5O1A8MbMT(_EAGV/.b153(f^DFRSV(G@L]dQR/B<1V9<[BGRd1R;[<\-I
]^A,FMPRQ_=f4T(Q:gcWB(A@(172,;:-93?Tc^75HUVON:^DH-^gTMPS>_3,Efa[
)R9Y2aIJ8(.7(E)Q#5_2,ISFD=V5P])G&-LKX&?,VJ6/^?P&d]5#<CK-K?W]QfIU
>Z@;_9[)f_\.,B]]#PO,9d[6MgdNA)J3S>b4(bV)H87Y<QRU8;1-U-9YVOGG?#M>
Ye==EJf-CO+[ICCNPM[+7Z(/=AXF?9QYOR;GJ(#B0RC?>R3_N#d.g7GCDSDH\INX
IWBeL#\(HDc/;CD>-L>Yc890a2N3#ND6E9IKPZ/(+gQL@R?F[#bIeJ,Y/:)?CN)B
D#0J4]AW?_8:<BIL;U6GId#-RZd;RX0T#?)af]4H4)60:_MY&LS[R;_YL\M1[,3U
J59^--:H:++@\Y3LQ>^_W0L;)QVN:Z3bK)8d(/3#\+GFHJZ1ABQ)_)7J=ZX;TJIT
.XDZ4MN]g&&,aRI_8aQ>ZW@GI&DZRRY.L&GY=#]@?bF[TcMa7(dCM\,>NbEL;_a?
6ddf=/&BD>857)D9HVA@</YYT+<4+\:D+cYZ67+BOZ]<V+e84Q_T]gAPd+db:(>E
.8ZRUX^O^JL4c;KT,;c>IUQP/L2-Sc6/#K;@F3g_YPF<D.V2\F(^48R;bP\M_HX?
c:]?H2VUE-5IGPC>32B5C9+41aLU94&=Q4Y@N7()X-)-.WDO_<GC]>NCR?)]@=2:
8+6aXM1XCPeTU<Ve3P^FJ+3J6#FP=gBA-SQde>/[V07>@eLGWU:UNHFK^>:7LS4V
SbQC^>9-02<Y4?Y9C;^aS=.-BYWT).5L^;P9eL/T?eQ7<ETRb>\(BX^O\4)T^AT^
Q3<7O]<AOT=(.CQN-)&1(I]:3C6d@<+&;-Y.Y9X,Y;A.KMIRETZGAQU1W?_S7.MC
^2>#^BCX&EA-4/6T9CEZ73?R-<FZFB925J]PKU)K2),/O?BD&eX\dM)P=9LU;J^5
NG;T22)5N?#/4]@X^6&NQ5+-U_bY4O><gS7=8g/6HaBdBRSY26>]/[64<:M><_dB
4@(>H4<Ma6KB>FH=>M?Hc?##1833b#8dVPDgMD9fD/39+-1N96>H=AHe2#GDgZ.;
G358C:YH[^a>d=R;[SaAgc0BBT-49g^JY&,)ZJX^3f;>DKW>;)27/0/8;48T_VO0
]G[@6GD;Y2ONbLA\K#5\X/@WKY]<,O(6V>NI=JO9GeR-@95YIb9ff4&bXc82Od4T
g6.C(<TIEAI,FI)L3^1V9=fIOJbE6B1/fQ1@YU2a=Ne@fKQV\FN79c/(332F70-B
#KNB-QL?DG3J\0>G#P<?ZCM^#8Z,9_M=6_Ba#fYAgDUWQ]:(/?V3O/EgO,R;?R);
Xa8:H_@TOcfK?8H._e)4M.2B)A](+HAc?XBLg-T-DB.0G5f\_5.JMU-@)J6X,/JL
</_R1ZLVbOT>F2=\d.(U<QN0dAJ?G\Mf@H1AL;94T,2.SN-6L6:.WTYT:D;a2:g8
^N\#G(8/feRGVBST<9R^85RQ6T1CX1\f,dIPDM[?DHKWJY9dXC+RB835@D-S7a0K
/[1RVb)ZD(:#MF(?A&CWa]-a9P-[,H]ON3NOa(T]N.J<_fVOHSg>J:d^KMT69SG(
UcJ.S4;+:1S:#2@WUPb>g+;^MAcHDc_FLUJ-NMQRV-(?=HeAS9]E.@VZZbX#6MOb
M6-OKDU80]RC)e_b\3@=4)Z:cW[C+.6G[Pe-N45Fga_\<R9YU2&HcG]P^&?-).>g
9FNa=C1)]E@fBW>=/&EA2=/&H\;g?fQ,1FJ5ZDF3,TFU8dJK&8SVSWCV:67Dg&eZ
c164@ZLX7/8X@FDe@T0+4W(79YHSe7Pd#YLI;O5)ae;<HB>9@1L/[G;=/;81)+WU
_&9F-7AMTI(DB8c#dcC0FNWQeKe9BZg7\/,/-d=8CZgc3.X0fRH(Xc?BaAF_=]6,
02a#Q)f\C)&3F)JH>TG8I8LO,TVf2<AbUXDD-QYb80_9;(E]g,@U5Mg#DMbBJV7c
3P4c#NY-V&QdbY3Xa[(_7)XUKgUN.YH-Fed05IK:JcN\=L)D\/2/a0_f6K6c]P=S
X0VO(02GeS[IQC@5ZFB21E;cIW+eJ9TNNS8LY0c6QXc0=FC(b:@Sc(^UBVd..=D3
Q54d6.V_fT(NaaOO>(^1:A)D[Oe\V7K^f@NJBIHUH_Y1MTN4c)#9JZ11DX]U0daN
_@MHN8\S3Bg=]C?H\g9K_K=V(MA[F:S&=a7LH?@e40\XTb@PJR5[8T2,?&,SJP2-
&S,f(IA94/5M5IDIBF1782cJ1/LB67g:\G7X/,XW;Le4=b8&:V_(PL,c372f=067
U-;Yg7JbG;[>&?EX.++Xb(6f4RaB02dV;N-XZ/22G9-X(dERIgE>U,T63G18[@<S
QGb(N.HD?-]:Ga+NRU^&(ZM084L59ga^3_Xf@B.MJ4WXcS#UL6MGdf/-I51520_F
9]IX>X2:>#K)VF?+VBd\N]])M_.UVOBRVRD/d?YNGO60HE@A&59FU<#\G,PW)[6]
M@QP.15P=^3e/9YYARWN^W@e#PFbA#UfIaF+.<_GK/I5636<KegW@FKeF9PW.JG\
O>#[2cFbUQ(+\F9=bCNC?EJJ5(L;(CdPQS.ZYNb47BVJG:JFB/8FSBJg<OfW)T,5
0CS<1W[/)DdQ>L\(Ge(C&19@<2H+,bLZ5geCT1Z.YfB\H+)Ja]g(.02UL1AE5=V\
2V=cc/e4XOBP.A91aL\&I.0+(OWJDP\27e989X<VObW_MSPG=P3aG^)^DKD]:9]Z
8@U>O0WJ53&BA6J8]9a,Rg:SW5V,EbA<&L=gV[A<dRfPA#0OBHE-PLGbZcY@<Ec<
fg+2Q\[),@c+5.E2QdGY&?>U6=.:0TgX2MW285JJVQ]a6+7-[GDJOHEP_#YH;1BI
Z7@S2/L)^gJ_@a5><cgGQ?VHg=?7&gEE(05TQ)3FZ4F<T[?LU&>9)@PSX7=7^a-f
Ua5P8<>cd/S<RaHS7N@aOB&6/KHC+;+8_G.c.K2KKd8/aUR?@.-9R3L.-32Q?84d
:Sa.QQ41/bHIE4T;I.HW.7ACFP&C\d5X11,Z.UYYg6e8?15#fM_]d]_0I@]O]<8U
ABab41aYJNS9EX3:)Y6/&cdU+F&[EEQ:&C8T3^J4L\0G1[I>2HU[BB/bG:0YJ?Q^
AN+FF6J<Q+6W3KOBD0]XC_db^IcKHLOS2G;I0fROB^OD9Q2PV(5@)dEHbVX]OVaY
H9YW3fA=9a]2H52GH39KACPHIAaNOa^SGIQ,9SEBTTGL(S,I<b(&Q[a7-7,BBGR+
e3N;GB44^fHdWe?H0_8FUUPV0MC/:4SDgF8Y&,c4XAd763ZY?E8N,NbH5;,2538-
=SEB+G8U:^YD&[g<Y;6[g9/1OEN8GbSK#a3VG;LVJBbPSZ&5OY1bS8H#Z]Q4+0C/
\^Y=SR<(0,QIVBFY9U>3?<H]-C##Og34]BEMIR:M,[PS;>FG9S(.d1S1<)2Q@6A>
H1d[748)b/Q6QKV=eC278N:>3E\7LX@K):45+993+9DENMY/USA.RfKM@(a5eC&1
A4E3a7Pg0_g<?)_V]378@C-Z3LTFK]5,Ad1__bB;+B[5\S5MP\e&f3YFcYc=T&Z#
E(6:E596CAVAa1.eF@RFGYM@&&+P5aX2CR^=9GE<05>dYc#dB)8fW>-g<Y>6]KM\
UB.&EVH^bW&Z8gY&eGCb>&1e^7-[X/E0:J?c(R)+#Gg<(5GF[G>4\OZ-MdI9J/:b
#I]1.=Sf12Y-;-_GRaAG+Y(MIb7M)dVSJL=:0bg6T<VX&aZeb<U+:>N]8F+?6;?4
dbK)WFX5H.59&[>fTfLA3[<O;9[(2<;^S.cCM4DE5+Y36&,X9[P_]&4Y6/6OSa5(
8J?LJY&a?VNC.0]:WW=RO?AB/PRK)(J1;g\BJ3OPb0>4&3I?B+++&;#)Xb<0E3@=
E0>V)RW_A_063GT^])@G>&?aT.4aP<1f]/g<YBM-QNab/>]8aDWN:Fg_NBPR\FT<
0,af]PFaHEAWR7ABF,a2DZ.dUUS(BeLFR6L93_AC@9?_@@OGgcKEXcKe+]LC>@#b
C3TH49D@/.=SHY_XdN\GO3c,)_[>Zc7LH@N?a97c@9bDBe3>G2TBDUbK7F-5=XD-
(cbV9=LF==J8M+QBcJ/BC>dUJ4KMb^XG&4Y3Da(G\@<\BC>\CcFW?fO7U3U(_PI[
J2IB=Q]EfY?]#F\;]?2;OWQ))3H7[2bF[UaK#3HW50^&?\L90^]UVI8-eTJaW[._
<[54.EIdJQG>8\N#+/?;1+]AO^Z+aNK-8FfWaN[YgW#gMQ7@W9eB@]e&7WfPLKf[
FcEFY(2#LG08+HK/)E/I@[L[c?JBYIFL]3,DJ>9-40GGTfY,=3;Nd5+A6OHJ>XPg
5.PA2=4HW8OeA0M+RINRORVYF,<MZT;01;25RV_TZH(eA&f0;?PMOO3NO2<Vb6^[
=7N-5A@_)dd>#Pc#8PAW^/c7fP)1)]f=0cY:F_HB,=@I2NcL<C3.O<#M2=BU5)bI
=Pd.9H)LOR>T-8@#R:,MXDN^U.^SP.a_3/\eT;O07/)HWA>eG7X^&0eLeTCT+9I&
Sa)ZQ1B@?HXIK+Ldb)?>BO#8Dc:+P_1c4]1g:/K#HD>IcV,_V(fP:NgULZA>cHJK
#OQ=Y])RG2T.]=]4:f<<]L_+>_PIF33.G</-LXT)8IcI&B7R?(N#69,[GC,GfX]>
,f4K;Gdf0MaH)CUNY\^:@a,=Y@CWA3_a,9NYNg?/07>a<X[.Qf64Z)ZP;Rd#-SbC
Z:=,Ma3;DD^)([aY<^cZ&SO@F5BU@S=KaILHaKJWMJR2I)__)3SIX]SFJScMNM+5
3M#XEFVSZ2:d/(/@O31\T0XOJ6;:Bd0NB+?:XU0\[F+H/99Lg]BIQg@3(_agcZ5U
\3_KYWG7e0,.,[(d45G^K01YaUQCXD^F[]WO^-KLN&=B)c0M,]X;c5Z\L(+BYeC:
+GNN\8;bB193(7)BDFS>BP36=+>L,O@PG?UEaXB\YW:\GZGN>0f](6)RI+N.11K\
FXJ)6)/==_OZ?I-]_\Kc#/Y&2HRI<ZXa:/V)[(]SOE3HZ5B)?YWeO4bRd,KfC^&)
-\_Le):Y\IJL.SJB=]I1V[bB1L5/&EACG(bX)ECD3b(VH(-I<3C&)6A><g040G3]
D+(-THb@82G9(P:TX>^^N\L?^5bJ<=2?7IUbQT,532&]KD?6Y^DUICJ(IHT,-[FE
Pg9G>0PXM#?cT=W#U)VGB1JgNRZN&N?AbNQ8Qg78FBTEZP-]_B>5S)FR_7.deHB<
R@5E4Yb=)e<]b,\[VIXAf=Q0U@0LC/LC,I\_42JQdG1+O=c@aCFC657QG5T^N\X)
47A,&cV=^@=T)M<d3EgS=(#Q_AHC5?.M&((X&PdAO3-3G<W81=LCK.?XU6:d,ZMU
9<5G52?/0O\E](TdU+EBDXCN0]UIN&S2fXdfT+AQ]@/_CJf+7K+KJ.dDFgOC4.@4
HObQ;4D6>&@M[S(@&N+I/S?&&E5g,a;d@K@0QO,FfRI&W;b]Y3fJBO/B^A0P]/\(
ca1@AF_1(?X3/08C-K:OceP@\BbD/ee1M3D;CYXa)2#E+)6IFcKf1Y+6;2gNLRNe
3Z4^.B1f5#/[]-:WHK\V?6XBR58A#Z8\b>PI>>FZZQd:JT&^P8),IUX[SK=F0P3C
+ER9a<3[WZ6a=We#R8V2@Y0/<C5DLQ1X@P.LUHQT4JgN]DX/PC[fUe91b1)e1<LJ
1M@D5e-)BL^6)-.XJ(8Ja5BZUTSBZN+FA8>>:[@8LKU,22^/CH/QZALJYN7>d(E:
6@D=bFYd^?N:0g+dX)21[Z5DTc8)B-P,;g(6>WNRP)6;EETMaPaOK96.EZa<=Q_D
^ZI\c+<&(IR7L(#9;YFQ53P)9U?d/-R=WVPN<T.GR#c6WJ?W&fDOQ[<4Wb^]:FTZ
8WII>:P)SY_FXa1J7^:f-508Z>#cJd[[(0@d<C<.9+478Q7U+fa[ceSd<KaK)/^N
ff.)HLZ1@71OKe@3VNK&MS[9YA]Ab=/dW9LV3a7dEJXB2@cU=7N2KC\(?VLO?DK/
H=[HG.ad?BK.5.5A^0Q[bERL9#eEYOD/75dY-#Z,a.P=O/T9E:Y7OfH=;C0JfdNe
EO?859@:EIQb-9#GYJO[]/?:/GP=ZKX\.)?C-Vd;N5;WJ>aaK[WYf(Z7>V2g1E@5
E8OD&g7aL@(L&e(7Bg8DaFKFJ1-WeaR3O+Z1G+>HD-d[E1@@(8W#<U3,_eT?4a_D
DP&GEX@C=&56f>LgN)Dg8Z.CWde[)dDG8HGG#I8e?bOTFX7UQ;@A8_,>Ccb^2f\L
EJI0IV.C&^gCZQR=(]9#cA/W2PH;6\EBQK&[_J]K\VPJTd2Hf4\43U(DT#UgRAfJ
>FX/Q,0WGFF5GYI[2,4\LEPec9g5;=Ad=G\J#g):f35W>#KKM##3RLc1]aW_7ec^
7<8V,(XdR+()G^B,XP4[eMXPReQ7gaNJ/VJE)F9NTV+Q<;\ECWM6<=]dUPV9\OMg
+=U:WEKSYGW.5D2-Adb0T3.F9#cd=0I)5[,1NSH,eFT8W2]a38:4fC0RL)MSeFQJ
R095@,W<_f[f4Z([bFK4OH_8P<YaLUgB+T8c+))-2X7VHXF<W,0N&6[DLU>D/fea
d.e3FQX\f[+8-]Q/>g@cJOR7[)LNH6.Ag@WHIIf8/0NFAB?;,c77;c][g.gH\<R#
J,+J][K6MMcgZQX+F0W^Fg91>aH4d42R75JWXJ-K#JgeQQBM[V]G)c[WU-AHB?13
2D<7UR\C8ZG192+[XFJ6(_EaFfQ71F^.VG][=--2Y(a.XR?@_MVd;+#U2N\2APF9
W,fUA+We^P_]>;^+c1U&T.NaeMQS2W2Ua_70_eMeB&8OBff;?[/[[:U@cCPZg6Xf
H+H)J4FRReA],SVf6-2=WTSMKH.J:KY()68_GXS2aQg_eXL@=+R1ZD/X8d(@aX4;
3UZ(J2&GTO3[JW8C+DZ\OG&C([+3:9)\)f912O5]K/I09H7#:-DOLfXNUfM88YW^
CDZ@AcT;\XbMLI_UL_/H1(d1-Q/MY_a.@L65M&fbf/7V0U=VUf_.OD>6H<G::83f
DPLScBS^RF:SQGY/=+dIW?][g;2&UU^AbNW+.gIQO2^X4/IbAS9f)IMIKN>,+O5Z
eN?CNR^[Qbd/#0(fQL<aC9@0;>?2M8&(WW?R-#SC0PSS1cAa@R&Z\XGG==F]=A2g
gYQI^[[PC0J9aY_WL.\J_VE;C,IO]9E?PafE[BXE)PW22?/@9;N@LDc&ITZM22#^
e\K#^KNF3LKc3c8d3J=B\B1S<DOPg9]QP>\3DJCe\\]@U\;Aa]&N25b)6M+,(G3:
90>YHGYGKJOSD=a;V&Z6.W\:eE8EVf6Z+/+>d<db9X?;eK_d##F83+VY5>7?3=?8
1##Dc8(-:;We2eIcNd,95PKO3#F38X,0X\R3JY::dF0XJ(F+2NNbQ(&WHAOOf&O0
^-3FYRW?PIYK#2+4dJJ_E,UHWeBbI>7YU#ZV)W;2;82c_b_.QP7S^+[,gLdJZ.K9
UK5:F0\C=WLQ9AJQceCP0e_J.e^@.H@U>V&,e/C23XgHGJG.4.ZU)=3OAN+I.1S4
O3d[YHBagBR/3)Q(/US@+B8.@G(SAXSdC0^JU+#gMBU2eBO3AYTOSAO;^>K9EI.X
<R#.]3]-\[eY]N+aL23@]Y8X]3(3&C][L)U]+;P?N?VI;10Q_f5B)HL8\X>H&:D6
_HKdgYa3YLaMQF[3Td#P(&=-@4+3:Z+e1SWCI>X5cTUPXE/__N6XC4NL82.,88),
CQ;2NB0GY-6E6]/ZTQU7.-+Q:)0A>6IH(4A6;fA/MQ1d\.T;\KA+;OETg(W4Ic]]
)+A1TB/1XHc]Hc?).--e5X#d1Ee8.BV^eI7V=A&:7-2@aO.PJQBR7fg<[#+WU:FR
HNS9Y>EO^9#f50)b=D/Q+Y:SQ7?\44R80,UT@T:F-6.Eb0UTB&ARR#YK7;-&S;Ce
Q:^UO18Mc,=JA2QU@c=UXZ/.AaJAYFC:K<QWS,G;;;Vb7DQ;c]CQUf4<1U4MXMeb
/56Kc=NB^P;B;9NLGdGS(J;.TD:@=)E[M#??TCO<P#d@<BT1O9<CU?3)P+AACQcc
4GFC:6<Q2\^gWT/023aFRXSaJNZ^G:a0M0<L2M(23&]:4AY,F,ZfAF3UG@2XMd=.
T,T&5e+Y^EMU;L>:59[X?]P[<>\J]Z##?Q1:b7KAUO]Y,4d\55GG\BG\M\0YG0e9
e3Y3:6eaXa8=[5eAVCNCJC&5&2NHMGA/NVA;Z6:W&)I(9]#M084;PRRZ5<RfH(U0
L+b?gU:AN[Q5]<H^ZG34UR?\LGM00WGf-e=<3X3]W0[67R:Qf.W#(HfTO:5R(O9]
ZQ29_T0f@TcCDUNM^[XI0)fAg&IDLP4L^\JbP3/fUL]URM-]QdQdf?7F0aCBCc&I
8OR[7gFeOeKCK);fVWERLDA<b[^C)8F^R/X>1ge0bR2ec2Y0VIYBS\[VNXG7\K:+
MIC8H4)DS_MC7ML8d_.@IN@O#RgPDU5fKB7^H/eYHVBV_9K]IZW8Pe+<OJe[@1P1
F<-43WZK2^\WFK7fL;P>b45^P0ec0fg)H_6CaQ<+0Z2;QDW@^DTC#:9Y>[4,\0&H
^T)B-a+@a\#F(VE,)DUg>fecT_9V_0&5bJZ<)_>#S\>S:W-UgO1I:b>KB6WX4GE4
)@1M=WRYe1b<eF?4b--6+M0MX^#_]9b+DY=EWYe,1SM2IT@]ed0,M<U4#7MU/VRK
)XG?5S^:37/@@<8aO))Y3/VW6KBYBa0,bU=R#N,P)8>0fFVa](010F:\;\)4;;ML
+)6CFg5g)Tg0eO5<S[NR,Sb+FIQD[0OQMB:A4f<OCG.GdcL53^bX\Fff9;)0]^[L
6Z;W+c9X,H<PG]Y]UBP:bT=^f)@?SUH[[ES24dL:1.SJ8>Uc=;/AJ9^c2BJ=KHEH
8;4\]59:-dG5f=4a66=F#R7;UY7L72fX[_),N&/(JR>/c7bV=d184;]YXT[T,+,F
E(DcFC87NB7gFMBUK:BaIENRM#DL[0B<Yd3;Ta9LDV(E0NXXXa^(H,c4L>&gS=5O
<X#8Y]\=/KW]Gd;@(>/1#d8],Mf7<[dM>2ZBUd&I5Z.G>.G^A.PcT@NO;(fbdC+V
g1ABHBV>>HRSU;RN8Q]U31P]gK#U^O70@(>ZE?YU7Pc2<V\=LOAOB?/Fg)UY^#O4
.+VRC5\=d^ZXY.7D:N6Z&OXW+8=]U9QC[#.?T,:)=Qc3g7ADQC))8d0YUN&P1bcS
8P\D]d1^OQQa[cCf>_WcbR_[6?[LX;U9JH+CY4Bde:XZ>dd;21[CRK8<2d-2CbET
OMBUPE.e9EJ4Y[dKY+3PaWScWE<@fNcZ9<M):C^I-JBE\TQV<-?OFCD0XXN#.&PL
><13T=c>5-5eaZ)HUSdcR.EKJEBE<Re&c<a?-5O+[:&YB.7VBN7bK:\cZgF7LTQ,
a?M+:EIT61DR#7(IIUdBU>[UaJ/?0E.adAfLfPVdE;H@N@E5ge_eMJHbI8-b6Y(R
b/\C.GV)Vb(-D<4:a54Y#0GCf_1:I[WaK&YV2IL6[34AL6&dBgL,.<9O9G?,-c&Q
=Q4abg2Y922S?GB-g/WWAL7I:[G-C7Y2^-cI\:P).LYc^][UFH&W0gQ9D-70BBdA
]0H6R]E@TQ[Y00:R?Y@fM5L(E-G30,J8#\f.(Q+5+8?8VR^HO@fT8]]SPN3(PcJb
7W>8c4DZ8@LG([5f8IH=).ZL--[#>+&beH.fMeACOd[C-b@L-)612VH[#H/+TNKb
<T7LC@-3,7UFWG@e872JACX9D](R4bIRABd(Vdd>9)CENPc4D>GYZ7HB/CHD.]#e
G&HU6:=S#V-BaEKP,PU_+TOR5-<PPHC.-CIA@L,&YSS^63\5F>Keb9LaBbP>^^S.
a2#;13R=HOg?I#:,g>IQgB_@7=]:KaD,^f+?=;/DUZG+H4UK&1eS)Y?+X5W5c>c_
I]+E-NH)UI#76eHe4SeXF11CDFUL9;RZ.^\c]-PO/6X15VJK7?AP6JWO[F/=]0+V
+NUX?^AbYM[G(A<1HdX@53(148;YV-C;g/SI8<#SB8SXW,@G<OEJ^[+=+gfdS1HO
0VP&=42I9KBHDbS/D+c8gQX>(fac#dZbMQ_4[f[E,[(;UC0\XT?^,;@:&.M9@T^G
d:YPH3gg4=?c882PHCONe=RJ9BYUP\9]M_K2VDP?>A+eT=#D;327+FgC_T/5WJRb
2_(0cDV9Y;@04[bC7f^D]NK1HgR8gT:G,F5[XN.->]5D-f>N#+OG:ea]-V0gR7@K
\POg3.7<_a2;MQ,D2O9V[C]AO:<?)=2W.B;1/YM1HNg#gE8R]bVcd?Z1b]L)5A7Z
Z8g89Dc-[Z3NDNG/.f.C[#2Fg.36Kf(E)D;2-PGC=PRX[3U#9_)J/8W<.RVM8N#+
9(C_<Y)\XI_#A)YAZC(2MS\P@eKO?A7=,X]6YZ2^M36dJ9R++cgS4UGAUgc3JeH?
9QJKd56J490&0(1S(2Ic4&A8OD;XB79eKH#OF;PA&5,[8ME35VeXdXK>X.R;V+P^
P7[M(@H>4g62gDI:dY_17FT/Z0HTIEIV)03LS7QUeA4?4GON7]^248fWZ1?X#D3f
]-5]QB^ZJ]?dPR,A.2.9D0J-FXM4E>^OY4198J&MIJ6JXbXM&[,,<fE,#a9/V7>V
Jae_MM84B]4<?@#OLO)d.(7Kg0;.&[VUeV4=QP>4bcOgYR+XOY5]+[bT2S2IN3E4
D,UL(T,4-f_K_HdYWe:TgGGYBQe2MW4VN&)Ye1H30\FPf.C=B\&I?f8b+^45<1@S
f2@;X2EF/g&47DQ+1M]8>9B(ZTTA?V=Y0.=+DI3T<#/9)(Da0U_A]+@[^PK[P8^C
e.G^W)3#SM41P#PfR#R&/4OYc_1_(&XPgI/_aA+</DL(T\=LU=<^_5E(/fAJ+YN4
dK=YO(7ID1KSZ2\YXW@03Zd5,28CYZY>gH>LAUfA:XZE,0F-^LaB/@PRH_D6IM&7
NJB1+[b5.OWaD#0.gGcUDG<W\\d7:_@#Y]#CJJY^O]X:Ig0VSRO4b,8<>Q.fOJHL
O9YH[0_0)Y^+C:RS<[.@c33gT\7W?5@;IaV^MX0MSYZFS;W64A=L41.MJ?NVaXU6
f3=U,4d;-=.=N_-I3^(D[XH172_gELR]__A17M19S);O\YI^)XWK(#I+(L1>]=5<
A^6RQ,a0MdeaN^&U(>M.O,a2;/T8)^69]IBW-:g7]NDG:1O+Sa4+fUQEA]=KP2ZV
e8._PC(MUJ&,@-,&RbUV&)7+34^;9M7-F5VTd0baOA_KOW-a;]\c,9WPNgK<XV@U
CJEGM(I7UGG;F#&CQ4a_T51=e#H:\M9Q1423S>#W#L=7-C#)/QYHMT]Pb7GXA2&\
PNY;LFBZW(&K@C7gYR4@=g?dS;XM^WI[5XQ5@\f@.L9,a53UEPNPT;]IL>P3:(7d
)I.)LaIg2D-B)a@EFBK17Q9-OB96-\I5;G,V?eHJaaV6]<AJ-bfe#6ZD4:L:TRQd
Q9BZKK<U&@Ne+,/UN3W]-DA&/^PQ;Q4J]H=GJW2@VERSfS-&>f&OLD/g(<@fJe&8
9=2SfH]_6P>N;fAe\D#0S?O0_A\OLQdJ2De6<GP(JZC-gF&YY<6^fNZE^3CIW#Z8
FZ.aA=Mb31[>W^g,GMGAQG-TX245gE1(Gd[93+F8#:4b<)<?@U+NcXJ(:g70;&,e
3H5GTbfLW,1CRS#>cR3Q3;V?8GeGZK[.I0>4aCE0U5_ZTf^ac1-]VCf5NI9?#O?.
9<W?QU0Z8C1Od#KUG3T)+U>WZ\:^15gKV/J7R>Aeg33d8/^IVZU@9e]0XPRTbGI<
Z<\@;gP[+S/d&2&_[R^CeWF<XM?V5c4+U(b.D/,^KW89)O>E,Y]+Y5882ASYG(Gg
NcEQ\8ZPDE)<Gb:[a/O1d-@S0ICg8O1N/28Ie>g3CMK,-[MXC.9fD.U/0f6J5=5A
FO<^+g<T/Q;KaSL-?(T(C[_#OD<<8+MJEPL#>URfB7)#\9(H\;R:bGH&9T-1S]FD
)b)gN6WBW+)FV]Sf\MfQb_d&S[MW;H27aQTa1BX0IcUB2_.af\;9MI.JU;PZLWO,
W^#J7Y28?8E&&J9C((Ld@B7Z>AWDGN8dJ=1&3HKU<[#66MC,,WeI7OI-gEJHJf2a
LVb5,F.Dc>MX\.URU8)/CXZ+1)-b39NB=_bU+<U^TN<U,^+]4cUSAfg;Y_dYb.\D
DcgB+UBgQ][P)g+7WD^C1,4/aQ=129NOLWUG\2Na5^2V+/YVfE79>_Y[7>W>;a,S
NK6015[[+HUJ5YJ1B7]VN78WMIaX<<70b3F<HM0;.^:K[#7G@\C,c:OaJIPXL2S^
Gg68)@DOgNgAc1/AG#.?LW5)C@e7BOR4e)d<7S_cY(]DS3cH^[4a]6c.^-Ub&Q@6
\URB8:C_9dHb7P.XW)JCN:cK3Q?O\<+N[28]+O.;bG);]?N1^S7f\&5/54Ig)X[P
UBI2Eg/F/()]=7LT5_.bNA^fOE9K);9(YP:V?e;,Y2AFF00TaCQ4N:O,AU.GWKF-
SGgC3;IR9aD3+C3T@.UTF6.;SRacM3&@Qa-V9aHDaXg^ISWEc+9-,_XG?6XdN[L6
AS=a/F;KOa/;>Y[IY<6\,4:bAgUf1(Bc=(O2[-VeCYf,b;gd.(-7HVEB2WOd;-QA
Y0T:<[2)PU64MT4[N9WRJE]:(RM,?1#Fb,1R1e1CW1^R8XP3)cMOY./2H.3T(G<\
/O.L>3a<ZAe+d+cD0=VIE7@>3Gc085.&U9V#X<^?>JJX53d)^eb/FgIH1\P#C)>PR$
`endprotected
endmodule
