`ifdef RTL
    `define CYCLE_TIME 20
    `define RTL_GATE
`elsif GATE
    `define CYCLE_TIME 20
    `define RTL_GATE
`elsif CHIP
    `define CYCLE_TIME 20
    `define CHIP_POST 
`elsif POST
    `define CYCLE_TIME 20
    `define CHIP_POST 
`endif


`ifdef FUNC
`define MAX_WAIT_READY_CYCLE 2000
`endif
`ifdef PERF
`define MAX_WAIT_READY_CYCLE 100000
`endif


`include "../00_TESTBED/MEM_MAP_define.v"
`include "../00_TESTBED/pseudo_DRAM_data.v"
`include "../00_TESTBED/pseudo_DRAM_inst.v"

module PATTERN
`protected
Ogb0NKK4C>b6=:,D2,OKV^O+b)R>fPD?RH7EN;7^6^TAWAEO6>[U1)71a8;Xe[0?
]#]J1^;L\9];Z[U()T;F(@P;Y/eS9\P;f2CY\;CTEA-)6-P6<V.Ag>\.SEXY8[DV
^:IJ-a#g0+N,[-/[#.134;cB0bTc:eD?-VFRGCg46@4A+X<>VF^^W+GUe]dC7)5Q
6gG<W+#&XUP3V=g/OPI@ICaQJ3MQ1H/[1g4U/W7VCXYP=5O8DT/8=JZ/O\=E]RdO
A;85ZBJg41&_\LAIb:O@0QS=,X\^F:Bd3&62>gZ=&aO9e7)fL[XG3W&0B[/S++>F
[2EaW07(c#<RRXfB+?F3/59b-,LfASKYa0e_DUaL:/4_f7b8I/L83<6.SdZ/7F(D
PRIPH#RfJCCLd@7f@^\0&7L]BW1.f^-^;22IgO)@0gc#,5H\Na&UZ4Y.GXTL.;=D
3:()&B8J&YXd_YG_ZbW^]J/,M.;DVB=<?@VS_8-e2f.F<gVD:EB)BS4<5N\-eNPL
<.]0R/+=+MZF+,N89g@E?:;+NfTe3Q-/8c6GQ#fBfL5:b^M_0RBFRJ:(\DO&E,(E
U-U9((KGTFZ4<_AZ7cN-)JE:<^K<^[O+eJUV-ac1?+9eWML=2-.Ugg=&3++[W=PL
H6=UH-@D/=3SSXb^+O>+N,QC-(=-#@-gI5cO93J-fA_9VTb4@B#JH?M,NdJK17_B
VJ;]Qf(8D/0A2&BA=Mb?9K?aW;R_7EGb0/V+E^IF>P(SbD?V]>(YOa^;fd\\<=WY
5>\]&Y0BZBB<TaaK.S8&;Td@)S7#7R80@W>Z5fE&,<d>BGLOR-.2)7G5<CJCDR6b
@9B-(I4YaF[.L\S-69R^A&HH8_]I1-FPfg1RJY1e#[R?7cY(^,R+6^-HP5W^5528
XGQK]/XUQ<2YS5gWP8OYUM07TDNC[=0>cK;g0I@[Z&MgODO)cL&+4,/2b#8H840&
FFNO#:8J]:I_&,,-fM5dgK1AV,[N1Yb:c/cM-DX/0XMd@CK<[8.#8E)-Q]241,N&
K51A_F=D(91bN;e[5&;J]89CJRgdL??2ggGYe_Sa/L\UcKZLFKD@b)79P[NK2O\K
2-DHeN9F293_K@6g]X&8eST.Pb4d3PWE&b/YF&B8(d8^e1?K39C[ecS:_[D1K4I]
5<1958@D:,W^cO5IHB+;81]@@TE5Q[;19BUcU@:PL8YCE\N5T9JV?@?0VP._T#T7
1+[ZUd[J]PLTaG@L?TXNV.52&&UUX[G2^O[<=X[7103C#+HE@7)T7YHJ5XN(RZM\
E7:\WY474KY;LNO8=2ZC1P^371B.e)cM^O9@ZD@;PNRdI_V/E\VJP>@TZ&Y-c,e7
_VBS:JJIY6QG:5Q4cXgELb#Tc@1-D\gI[H7N3X((TJM4#Na\1Zb@Z2[.gIVY_:Ha
+3B#DPTOf[2ON@Rbe8@2)b#BA4VB((XIW@d@O8#YAPFT6gM7e(,UB_/AS_]H-+E&
eA6E6[6CcP#YeU;2>0;BY&1RG9S]]<@Yd/WT?HFDF.3gD7Z]F2P4-QTVFf\PGNK=
BefE#_BS@JT2Z)4YQ.4B00_EBZS:8OOJ3#Q7gK4b2e<76PK,]g#W^\[<E)?2MBAF
Tf>bWU),)9,eJ<Zc(7JC<6bNd8d8_BaE@g()&gSV4G0cdc<C9\SQV?g/X=[0X</?
KF@T^>HT.\_ST]gd>R23G6[VHIJYHN9/33T(M)+4(6Kf^/4FWQ-2QR2,6EKD6SSH
)2cL_0U4SSQ243MbEDd4W>fA:52@9;E;@Ia#]QP4f])HfbaOIV80D\Q<XUDNXU_/
U97-gX/G&LO_J:\-LXgXOYPZG[XBMcd-6KBDE)BX;TSOJJeV7XCR:(Xc5@+JG_K6
WQ\eZNES-=)3#HPW_2?@d0VK02&^gCOIQ+#0:@3d[\C.#S1KeVO]PX(@bE/F9@cW
8BC_[0>86JI;g[9L4+I6/e;DI@7^4f\&e-1Q(TVHRg&WAP_&a+fV\3I@<b#F.M;a
TE9=MHN>b/5=Bb:SGZ]>#B+POS8RS_,K0ga,cFZa30BeG)8,KXD+\Md]A7a#LM=K
D&K-OWRE_N859M;gb>]UgAaFS@SV6dcJM3Fb)7d/+W.U:_V-]gS0]N2NO,NHQ:A&
YC\=4A:eD4M=[7#7V;L(:daZFG37HQf^#N<;JTQ,W(44@]2/KHDQA&1cFW_0-UA?
6_ND;4>.aY#DX0OBQ9VADT<9A<.@[bdg06]?=#>K1e/7]\3B_[1OSW[\PHE&a60^
&>PHW3D/_MZ3Fb8\_L,X&+bT90=UcRMZ7;636,gg=,][-OE2=0L24Ba]d^CSQH<4
FPY;B:S/8eJN\V4;K+^&W#FKA27DZP2ETS_+MV@Ia([P3_\)a8S[&a^C@\-Md,4<
FMNC:D9.9/.H;?EDd^E>,=G1NaOXfE[CEK-UCPE<R;1@DZCTMQ:Zc3dMW2?M^=+I
TFHN=YI9]?N6:d,4,XOQ>B/aY52dfe@;8GdM(ROLVH_IL\gaKedGGKBEZ/A0W(.f
.CT;4>_@^]TRGWII?L#2]Ca>,Z]O176G;<@SSI0Y6[>6H1UC(VF:&Y1f]5[V50\U
<7:(E;&F;eGHc?]RB9VZL0KG;+]ECJ>5?,T;?19KeK<f^S>QN3>)S3VQ:1]E0Z+2
TM#I#GKdSO6(AG>aHRC2CD1;4/?0;RXb#78SAf:@+Ad8;^;/(IKe^cDGV+c0HG2H
/DdG9_.Z;c-TS8@U-O]F,<KIZ,7[;OH2fHF2,>8cC4W>K4>I57>/9c/L0,f0];?&
Z+/=U5\_\J(I(,==5RG8UDT5WOD9gQaYL<abSE&V11dS;?:2_]UAe1cFZQA-^b;c
e9N(H0UdS3M0^^Yc@>N.F?;CH.HGS1UMgW6NR83C0=Z@?Ob_7#=YWA+89eJ4C/2L
/WF@N24gWGWg4_^f>31]4U-MJ>F[B:<bA_=K?/91gV,PMVS3XLY,^HfF2+b_VB8S
OBZWRd9dOCg7IGd5NIT(F)5M[FMLfW6LcIdULdDHbP@MWgN;a#?3T/F[W0I<=EfW
N?CeeB57>IXG),Y[R7S&DOE^O4RbWHa&OIDW]DOR?X3E9T:Q8d)EEG@3>:,H/#3B
TY0;C^1L_.BH?M25L)[CT)[SX4Z,9;]f1XE7-QS&7[c],,UGb[)M4P3>Y&DeJKBW
DF3aZ;P42W=N/W,MRCaW_BFIMQ-;^<AfF[T;H_KICd+19bA,bM@N628:3<SB+-c@
QUEd<4N^R.-]-S^faf:+/cI]5>@B?4_M:fDKHK)^,7GXY=C5?faYHgI#<86V:.Qe
6/]K.B+-QAT;beB=&8f7;,G:L8>JHXF63D,=.Z48NeJ?YZ;IM(?NKg75K/G<IXGG
2(IY.CYGH48H072W1T\<-]#4MH?3PC_>JS.LO_@2@C,0K#LK^cW&F(gQ-F:aT:O&
4NKQMV2Jf=#b)CH^H:/^7+X5X9?:TCS<QBRRZ-_.PD\S__OZCH^:CLQL5\^L@Qc7
NB(2;FBG9EE65@5YI,M-AENcEB5fKc7DcR3=ZW5B=d<5\Q03@-]EUENP_JRbZgPE
,/5/f7N^3NXIE?]0e]Y>2:O?8C)3J@=:Q2<F-/H@>d+LdE5;TdRWfC]5O4()W9e)
J,KZ_,BJ8)8Q/a>EU\1N/)80Ua:26If:LNeS<H.8K_S9Sg+W5FAM0V(:BcQQA.6Z
7O9V+AJNRR/TIB1K)2FZI@V7deXW11Y>;Z;UO:(6^H0H&-5eYA8+f^Ub2=?BMC/V
Gb1\;>dH((?-XCaI,N-,RAL--^R[9)WJSSMBVTJHZ])H,09>PR;gNf6)c(4#IdaC
e()ZU#X>FK8/8Ba(;TF5fX_WNF^DZ?JVQ^C]:D]f-U,FQ)(LIA8<;.+8d6b9\RM6
G>-a_8UG_=fB2+;gA^>BOL31QFQ/0.NG&5SW#5I>?:#5IQ,STe?Xd70CCEP7O5DJ
8FS1)KdOXd@aY57b4@Abe,:?I3AL6U?18OPE/dd_:a//3Q[W<ZZb5-01(S\)KaFJ
F+\RaTg#f&_]f/@\UT1eFc_6aGJ+eNT.4e2YLO_JYdZE_&.Xd=Nd0T&8./1P2P>O
8Z-ZZIV1,56]E.PZCI??VAHJB\FFW5L#(eBbF:4?_]ffYZc(#36Q9(NT+0KaEP7S
@G.3a5)6IO?=OV&YM/#.4ZQ)Gdf(/K#7)N#0@SR?S=77\e&8;1[<=PI3J7cH9]B[
9S3THd5(X_A+Q2B5fgLG@Og0a8bgDd2?[?,QbaG_Nb=ND9CT0M?5MXS3SgG,>cCD
#Od@g&af#@I:Y?/SG<0I^T.UMB#dR6U6@@&XN]4AT,=g+-?+c:-KJBQOTdUO[^+d
[)e#MB&QOf^f]55CV#PD3UXH55MPBU8Z[FY\WgGO)R&15PKff0IX2:Uf[==GPfE-
)_52eC,0&_f^e(BeKdS/T+gd>[NI39PgRWRYX-PW(3dc/SCBgO^=cC5fH4X4g;VT
)gX;Nd+fG.^W:,-D:eM?C,;=S6X,>dR43Of;FT9=,aY>a]-2JDc1-(A^^HXXd.#6
2>/3]PVZ[56UGIJ06ZM_AUDH/UBK.\cUYad:KAWEOLC30IXd56A^Z<B<Y&+^@Nc6
L@QIL6(7eXR]JFfY0KSd7J)AWgf=37[)<@NC;:dBA8=M&4Q7:K((C5VPeg&XA9Q_
e86cCd=>geYB&bLE<?N9^S3V<GY^HBW8HQ9\.:P68b7L0+M)C_,-cDPd[K32@UBa
ZRd#Zf<+()SZ^&fga/+-/T1VL59G>URC7=GdI=cC6XQ&7X2Od@C/]d4cEGR)<Y3M
;a:)QXVYLVW^;QcK)\FG(:^/YCQC-P01EEB?8R^0SgU=YK?D+,=\bB55L6+BOS8T
P^dKVVV10\Z^[.=4)e@/S)\&KA,?JV?U]Aa9eY:GG3#5d>Vb<4\HFM_VPNdUWSLZ
FGL#aKW//HEK992S9G]#BA@]2_96KOK7N4>c(F5P<]\AZSC^Z1d\f3?EB7^GL6.=
f+IY6((9+GH1&&9H@UY,?:H@2QgfXcNNKDZO,g;;3fcE#ET+IU@P1)0ERbS5BPU)
(a<18eeL:FFF9J&Eb<XM5A&A8P\H/G_A/O[gH8Q?)N(QGMb<cIP^6EH1G-)7ca_;
4bU12RFgCPeW36@1>?>c2e4WT3Z:-[(MH9FGI2::=).EJgfGLI>7F=[Sd0.Z?#<\
;RP<;e4f,Q?</Dc=H))Y3^a=3,S+f;LVPGI+\ZAXd?\BcY8]g#MAb_fV.,:,F6aL
VCL/VH[b5IK52=GeIUM:aE3)6b-8^#N=5g;de;ATN-C#0:>&U8TT[b36?Rg+6SZR
Y;5QOOe,SN+[H+R1SZ8C\8:4[(KG0?W\^#XBBB,VC0Eb.3X(YO554:T@C^f_[@8(
LU;@NZ#+/<>=E_a4P><45TJ=L=bI>T6cCP;@)2?)370S[KR]0=gJ>PJ^]#dWTWN3
f-&BM,dd@bPbG=6J\DD6S:73/b7c(A8D09:\MS]W&?T?BV-#R&g5QUVE2]aK^QP8
?C8P1#ZKA]L=/&aQW1<XJ)-cQPP@\=+]Q<@+3DRM3LY/7(>a\]Fg]_[dg.DKXY1G
V^NQKXb)G94#S1GRNBc+L0T\)WA/<DZVV0dZR,Z]7dONf>3<4].(45NI?@1=XZW?
=<KBcW3(Q/db@6gg#E6O/@1gJK/C]4;FW4CHYP7FULMGT1HPR>7>A64TOfS7JgJG
<KRR^a5\eA[cARG;Ha_SfJR8Ub;HPfZO\;=.325Cfe@(-3(>J1:FgNT:fVT=JKDI
4,K@PHdM=;T-c()E:g7J.6UPbBU3:]TPG>c:Y\VD5(1M[3+5^P-<Gd9Z=Hc-JXF[
#geM6TG(:,9;a=PYM9F3IW7.K/5->JeRJCTVLB+A[DH9GH]=C0HD3;^VaV^ecQH^
E5e\B&>0K2b0C)P:GHV+,&U1dbI,A10&f2g;,841,dVgO5cf3O]^>7?UcCS/W4@Q
Zc\4e+b@Tg4(1PXC28B?V4K2cF)K7#5g7TBB[GF@\7I81,OC&DF4923HFDUJD19T
eYBR>\e0VJDe[)Y5cD,BJXH+d)K.3E6W4(dR6A#66J<IG>QJ5:E<VO[;>=&3-O03
>Vb\>a8XB1LbAI^L0ee8dS\V74AEbO;5L_D5.HENR@.:/D@0Ff/-Fd401A-9HSeL
KH/Q>Y2?gZSO/D^1LO=TaKP.F;e8SJ>g+>SBI.dB[A)0JE7Zd^?6AZR-I\4NS^=)
Z6VE&W&#6;d/<C2K8@@@GQdgE<XVZVa-3:._&;.5J1PVXaNcf0Lfg7?GSCCZf?H>
V2WO-Z=e)G?63AFGcM]2X>>c3KC_9g26XL-IXKN)6U_R(;>Z?18_4&VOGVE?,/5G
&;4LT[f6)L1d0IZ;P@gWQUK.b(>EPAF(?Z#YNZF46\URXM.H213JcU17X<aeJ;aC
bU_CdMW,fZG63]\VEEP>7Z,0]=<KQJ>e&01e1TXO]/[b3A3)b&d\+>\9T[?HA#5;
Z10355RR4M(DB]NDY4U<GSUf.+31Q([,L;_bXbJOBP)C.Q]Q@&5RdGaO3+Meb6<2
3\K)I-J7Z?^.T_/82bZc:9=?((9[M02>IF[X7L8f7b#W+VeS7^ddL\]>[,UUcUI0
72/+G=O1@T5JE4&5fPYb<)/,ZFLf-G?b2be3Wg:-K4MEbFC:S(\Q@0IY583dLCD#
+_U1JME]PSM;)FNX#)^)/H<?cL#P[Va:@TM=^MF5@CRJ2cK^Q0eCRB9MSa5B;1L,
DS:fY&QJGY&7BQ/\QA<2V\(=T:5(e?8-544cb/YMH(:)-.+W(S4b]aCF,#+^^;Ma
,;&^MC_XB,V@L([BS=6G#BFb<L++0[2+G^B7^GZ(&cPcWBOLfN+7C)OB<F.@E_CF
.FaLAaD;[M.fUa_KUedF>>^<3QfCYIF_487W+eM+N@&26cL)+OA9#<;NN30U>\35
<:##2E+bC?\bLLXeda+#DL&YD^]^3Z#Wb9:XS;e@@fR[cHW.Q&d<,W,.K\]S7;DY
QKLKA^X/35d<M?f<WO_3UJYVdG9(:?UIb1^[1_d[D_+Yg3VfWBA@H41([3cC>RcA
d,If[?;C[Y6GO<_JZ:78c##_2Z(Ee+N#cTE#F48:+<491GN80;Ma[JUUHa74,W/-
^,^=ALK362T@&^[M6D.UL>cS;7.1U5\PH0g19RK73/QAW.e2021cPCJ8&e6RA&QE
2R+J;(H0_.>7;24U>THWI?/VTbFI[IA/?1@W9T<S_c^+[Da5GG45455,-WKU8UCB
,9b5&>WBfcOU-GD]1+HIRB.C6HY#/IR5/V(AfIB3RK/CZT6<VGJ@/3Y@^E?4cZ/3
e;ZLST^Og?2.IN>=2<>\=8R48DV^/GJd<f+^/a4(0A=/g9>/FI2WOO9TU04/8\;Z
Rf2Z,D=e=OBc4EAWeR6Y#U;bY:1[ZY;cO/^/U4ga_d^;6/B0(Sga>\R+,+-e7ZJ&
_&<-ZCN,2F2-&DPARS-Y>/S4W#&C[1aGKE<B+97e2SS><26&D,IH3D&Q.DQ:H?W7
67]KCZEB\Bc;28d+G1WH8#ZcUQIUO1#6+I_]GBQPW=eZXId]aY#e47T;T@<+X6HW
(WH2;RALa_9CYCVY;P<dZ-fJ[a<N>UC#A:[:-:1NKTEb?BHR/T\;X8(^3B821.MA
MG+A@A@V-E7OEI16f<H(V1_OZR;K/@Fc\[LVGOHMOE>N^Wd8\1983]KUb3<+SH(4
:1#9@VJ&AZ]O7>HXI5b.S.,K:U&bKIf1KEF29fUV+FMZTA6,L>8aV;cJeQ#\5\H#
(>5?4YbOH@X/a-7G+(3_fX>EN(A>5MS=W#LI@GUQE?dO/S\6A;cd,AL&XUA6&N2Z
_>bR/8L&>AW7Pa&=2+e30>6Gb[VY@M7a;H\_b8Q#XP8JEX\8@P3FE8#QcGW]>A@7
E8HYM@OA_g]e>N&eVN2gW86CZC#WQe/C&<OLSN1K4e/E)D[I?M1L;6/@7R^?I_Xa
UKV:8YZ?U<>&\5/ZI1b5&IWS&6>60,I&>0@U,?J,6R5OY/,+[,B3RJY2>?SfFJ\V
fWK\#/MNR^e3+E@]ZG+7KAM?9I6=?(D#+T>X6b\g/VM@(bGN+.d8JP0[b.(]WAH=
&P]\JW6G=)P1_DaP+(cP)O:V_fS[G=RHTHV=&IN>Ug6H3=VcBPLE5WOf9,WU=BHM
+S5QQ.Z5GB_6B0H-NIF8Z-_>=0VfK57QWba6BV4;g)7V>?AeV)HC26_a5E@O9\-L
_AEA^XWU^^R3Y68QS()LY9[@<ZF\0>fT,[KEfg/Z#6Q<Gc9]efA6D_0_<1J0&D/V
F7AbEK4dB[ZO1YeTFKb^_2NIdEQQb2>SO-a\7F7DI=SAP8X_Fg#AHOK/I3<#A@N<
#33K5@&BH3NcE-8>a4[G6R\e,]_#]3[37(G;@Ee^+Jd9?Zfe2QM8:,O5b?OMP.Z.
9262V)P>]GdMJ7,;]+/9:AJ,b[9d9a^9]bLb[Ub368R?3E0F1VC&8fA+\)/eK3^K
C]_0eM(S0]N]Y-9B+&]Ha3G_+DY+-SI9N+?M#90CK178;H[.B6QA=N^,.WOH=XXW
cUHd_F(V^867b)RYRX9d),=IR1(#>fWKEEUX5[/QU(8gHU)Fc9C/1Ae2Q6Me^Q+:
].T(@MJS(&/@/ODV3E,[5VbM_R37@4).8[0HXSA1a(Yg(?#FK+/CHH<--?7,_@N[
Kbcg+TYgc3T#M([:fUS[5Gg:9SEb(^<.5Q?#ZeS,Y.71d8O<cCdY5@#TcLB,Y;63
>/c\IDLe1QFVeQD.;\8Q4=Q:@4H,a#d^;8B94,F)Ifbe#fgc<3&(41\@eLE53Fe)
I;D9B0H7:cOLQYb80\N5dI=D7WZC23^fJMB;+THO?M0d(bXOa@=E7::^._YTdH0;
DUSdL[+EZRX4NDF>V.e-Ccg/7=)Jb6ePJ)/(e\K6Q35JP58[JKd@Y3e>#^^N5.(,
c3R&+E7._G3940N#:N_IN]JXLK-5LLRc:b.3K#Y8>2_cdW0/\=R\1ZaOY2_RUgR5
X8)f(TOO5S<-#B>cQ:2:cg<P6)ZH(IF@>f<[R):N>L]bA,M[HNeP_Q_351H8NP(I
GU5\=FBEYMW8WSU7R1_IF\^WWLX?FB+X?WcC8NWORPNXda@[T(&9K[RYFW-,-V.C
a#7dLOTJ\&eM9MRHU5@#_8RENF>5_dA7W)LfG;G0O:>J9R>[E=b3<XJad)B:\5OG
aS<8cIV@1EH>.-=7[d6U+->K5TE\fc6Y<?,SXGdF+1b-c_O\J,90(&BF-e;d:eO9
R11I8=/e(,&92==cHG>AY#2&V7-f]Y(Nf[2]4AO#MF6fVEbW_IU(U8,[@=bMQZSD
+/E<#?ER^TRIHTW<Bd/\^K(Df4(71T,34P&M8:aQ^7I.O\,-cg9AHDf@QU8+,Yc9
_c1J,8&?0]?<U8eQ^ML4Z_<8&IWL&KD3+QMg-RJg\[&;7]c7E\.W]O_O,&V6<D#D
<4371TY^f83S=/]fgRNSdF6[4CgI1HBQedTC<&2cC>?4LW[QH?O^>1M[V7?8[WD^
/WJJAOc)7SBW0HJL/9-U=449;QFP-6K9G=aWGdUM,CB&AAO-C)N=&I;M,e]&J2CT
?/d>U)Kd3N/N[BeOA]T:G(I<X0=\@Z+WU4;3#N.>5B3@9D;[[b#dG]cD^CIbAOMg
&/S;C:SCbe@KQGVU-F)N4+7>b:T7IScFG0Q9+ITAb/.24bJGd8d(fe0#<HI(1;0R
:XSb[-CE4Kf1<9)(fZX5a3S?K[_6\I?SGPZBEAdKF>#K7DDUdMf_8^T45ECdJgUC
>_Q&LALfQ_PLC(JT5E(HdQ(OYQ529[+),TUI]1]g^L5b1V^\Ze<TSYH.^YB3_DF0
]ZEE95SfM>BC[cBRcg52ADTIAfM(GT(LIHZ&I6A_QRBN90H0+#9))/dU74c=gSf8
&J)>(_J-SZ5=B970Xb6:6VX<+3FI)+LA:CM,A.H&\P&._Q?EC@_Gd&^Y4/.]M]X5
F=0?0HHZA5V@;Z[ZW2eZ2IZ(e]bC3MPa5Q0N+])0)RX>/_N<\&A)W,JBTQ,U;NEY
9d,>BdN0a#>f:d871S/XX<KTQ?P>ZNW24E&2L15W5K&[KfGH0aNEC4I_KPA(29N@
FM\K>-2_Yg5-8\.T&aVF7U_gAL+&FMC/<W<2P?24a#NI7D6+M+d4QG8)ZFJMfa+Z
QbI.S9a,MW^.0?9BPU<=B7NcXNTV>1[FCS(S13>G\NRA58W/R6&b3:dQVUI,F8:?
be_FMKIU-HU4P_.?1G((#X^X;XJ+_F/#D0:;5eQ93C<dD+V9NL:0D39A8V\F+J90
[<:;g7=#db>67?=V0dBdXA#\PMCb2a-0@]TbJQeWa9/@6F2]:7Z>]S]PKTU&>eg_
NTZd5]_^7>M\2?=G&RYYURHY.c.PT<#GFZRRA\dIC79<c]_J:O77&1X3^c^g,#0D
)aGQXg\2P)JdF]7832S1<=9+Z0VVU#&S/].<JF1G<(A-(fQL_)+HY[#](bdM+5]U
9OHINW3(4A/Pd\-Q^=+[ZY&61GY<MR@+[;[Z:\FD4)NB@^(YV1Q-42a2FCP:f_Q3
RL#P++c+;?=D+9\:bg[W2GJVAL&\a#b[AP0:,^/E:Z#+U94Y.2:PJJI:Y]=GT/)#
3Z2F0X_Dbd#),8],b^,CY:,6UNDD-15TK9Z/-44g?IO]NI]KBPdFOU9U/)Ng2_G+
/d?I0DPQJE>OA,B2H\[OWJea2T((UIRG=eE<COAgTX:G_KU9\7A)fD1f-RHY]:2:
Z;-Sd+e]^R)57f?7DOREOYKaGaXGOPgNREM<PD[+BJ?2GWE>#TfT9d?VYE(0>I]R
/gARBQ<FF2IVFBC&gT8NIGKd?IO@68gcSK+BaI#EHO<fI4:L6af:Wbd4F1.VYZ]R
E&\9a+PZe3?TgP,W)1efV32A-U-b0X1.Cc5F5T<:?>(2GUaII;Z2N]VDe)4U01S5
EfeOOULD)&,(;W=f1WIIOP]a1@eO4_(&JGZ#J^_J^WKd700CN)6#>Q_5,0=8XQ];
dR6O_[MJ-F04b6TS.B3G+bM\_W0462>/W4bR@#3M&XV2<IER,a2O++ZGgH,cXf^:
J#7HCB7A)=R)eDg?cW,:aH-MTH+_++UMB:CK&M,W&I1U;0WUFT2_,3[3:<\H92+\
I#YbOIN-\QH.1c^:0M9+:5X\TXff<IG/XO&2B0?g_?O0/(OCM:[SZ[O:?E]TCP+Q
.-^X@@>26-=b5&E7Lb];6R,FJW-:YJFVR\D#(Q^.-?0B@gBQSV3H=G-,2.-UgH(9
@V&^T?-1/aGZUE=f;]FML(fZYg0MC>PZOKOK.ORB6KHKV(@Y-J1<D[HK:5fS,1/Q
f5PNPK76:.ODE,cK2@IS4fWJ&F0D)35JY=2RE,[Na9HIKHc^=c=TM)@0\^V?Sf?O
.cbPJ9(?OgS2X\JJ2BJ-7T?cN&GFI;Pc,80bY^[aS[g>bCD1Me)+MPYTcW/Z>AW?
G#3(;]\(6?T-a9@NF2&PD8_897^IOUVB)\7U+6T^=bbO7)M451;P)0O<DO]@YM7N
f=@PR_]YZ3P6>IAK2a\&JEU/&Hgg??47T&4Cg)8PB&8V46(8RCVCN-K9STP?b9cW
341b]:8>2aTW+b;,K<d9H:C]R?V]DdWJ2\3Z2\.^O4ZAD61I\g82=<Ze[Og0(^:)
DOd=@6faaVF[D4FIPSL8])LUXD,+.[5>E8@^)MWZX?SFcb]JAYZ;Ya6A=:-cIXE9
gP)0Zd5(KOUFBS(QUHc4Z)4-?d1W0LE,Ve\NH/=L+TB-K>;f[TPEJRVO07U#ZC9S
GB9/\>85^HgTB=+MgRVQ&E8JLf00<+ZOP/:DGZ)a8S-_1,WDUOO77L<4b_/[gFL_
[FGG1QQ?ZdRR.bW,5:LM1MO0GNTa,JC7W&07C+F#2:U@[+N6JI(gEXPa(8>0=+HE
0GH+0R@&55?8^,MbMV&2,8^]MWJNdL+Ae9,+7NNM)e#1PJ<J&PL?@W7\<\Y;@)Q+
0C-GO?>=WNa8e+8C-C/N-cPL[G90<B1aYBZ9BXO3<]&=fPOC>V;F&O/XK_V8UW/>
(9>];e\;FUZNeI;?-[VA>]3_FEX70V4=c3WD+IC:F1YH[Nc.LB(DaVXQ<#D4>HNY
J.c^Y#Ed+OR(1;?=@<bTeXNJ-,CQ7M;;J:0?2(N9/1;09aaB_V.:Q+FaNAg_F]RX
7ECJ8dM6R8SK>/(Y58?MCAVIaU5^R-/AP22+\^I>-DNF\ed?8fAWY#EaAHB86O97
(Wd8P4f8SFSRSUHaCHBg?O_6;@_1NR(F8QfYJEH4U3=?MS=d,H6g\:GVS1d^PTa]
L2ME.0(@<QY^L50J6Ya&M:?.6F=R1DXeMM_RBgZSd/2Uc1AFBcfG7DNG;8.eMJeB
\c0M3C;e,d=DM^5VRJ?d#\L\UPV7(,aKFKSQ<3WBb[gQ\6Je,L7@],d<,0A-LDfK
MDW=c.TH9+g2T=?#V18PYI@-Ic1-./I/IQXEAULc@VPHP98+WFf6/<2d.3U0c]Hg
N#<LK(HdO/E)S[TQ2M/K(<Qc;_D-R<(;a/aM.OA@a2cZ8dY+fe<eVb(L:AU42N5H
8ZTcK:,+LZXR:Kb4I9J5@M1@@RD\:J?OR=9O7[GWWZfb,/A&XWMWD5\:-b_:^5>e
<VD6Mf.4OYQ\(^KgD3SFfT(F0G7HB1EFINLR2c&Q<Tg(Z.+0aUN8VV#Z&(50A6;)
:ZZ5N>KGC:X+G+@#FFgU\]JcL23NMI8^^\^gP\@?F9P?@-:78ZRBNG9g9:V,YCBN
^3aNOYNS7NLgVd,S7.&@)TG?N4Z:daI+>&=2W]Qg.MDP5:NR;eLe&RKe>GS;F9W+
Yc6c?R/I6EO^<gS2NPegcW3?&4d,]T#3NW&^(.6N-8RdB8:11B4Ue+NOR_4[]E^A
0D82Ke-Z,C45?F)\bZ^/16(PD?95EgfC\.VJV\9@EaH9G?gGcPJ/+SF0bL/V@Q)/
#-/6(MUO(ZK6XTRgb#6(>G9TZ[.-.F#DN@W7WeLS+MR-BI@0f\V9HU13;Hc.6TD-
E6/1:<.P7JTd]1+.E9;_&TEV0&dd6LAb\e22/[0e2)<3d\E5[B+7?0:f5/N0b(d;
NS\@QdIYKEZ_D]?]AL=(\/MN[/0QE\7\<\/0XQP1+<H:?LUEUK9dMLHcBMR0f>&O
<A4KVF1YXKbCPG2Aa,98J6_+Y#)-^H;F-0R-<^gHDbO&:bX;JC7#)UN<G&056e>^
U@2JA22X#,e]=OgU,=e(V8b-^<&N9VD\X+A5./f.4QK2YB3fU,)Yd94:JDc3c0/K
\],EcTLcXfb>KL#0ZN<:,:.Q=<,T:gfH5W.0J@RS?6^\,ccZI55c3IKdD0XA3I()
>]IUbESJ2+V\A(bQSUbW-_RWH3KNJc\Z9B=>5c:F)e=V_84+b^9\]f<5XY@CR)8=
2<>gGI23W@9-^VWOafFV\4UG@1OBc82cVZ0XGX>3Y<M1D^#]W8QDMBV:PZNQQAH-
Ud7TP3b^X&;&3d#9V98;L0DeP11-?UC(?>5;]&0L#)gHIW[1A5KaA.IIgOT\UO&I
dCPPHRZWIOY;::PNGA^8]GPAT6Z./Wadf06KLa^6(aPIT7ZY&5<2UZ=gN4:0O2b@
I1G+)H.7?:[JMV\G^)J=(6SPTgUSA=:_8[@CLF02YNGFg68Mc@M3R1TVXLS+;g_5
V.#d9L(3W9[Y3?XOKZM<a,1D5YbFL)d)M8c&:6dU),[=H\aNbSe#<Ge1DOFOMEU]
g9@&Y\_O_UPN&Ee>#X8Q;DJ@GMF/1.+5I.:a6^7>FLAI:(K0+,\KIW.McBaN(WX8
V6V8[_+IC.FYHeM3WWaY6ZCFO_;1+5c4X-=;Y84AQFLdHZGP1ETP+2SFAPDD@P.C
QGc6GIB2,X_./OSNT;7g+FAd>WC5)Ke8+GV.Z=UFXYA-;1HR7ga7H#XR-<IMfgDW
M&cH^]+Gg=#8fY_a=^&bZW[)GMWS[XV.56DNMVKbD=][Q&QY\_.NgE\)X;dbOP,b
M--X]_(7D=/(?W9IJ3cR].=9Z=DC]NK@WXAb0L.VCE=(c\6#\ZI[Q-H.LE\S]C(V
?<&bL-ET@fTJ;FXg>Y8J>-B5@/^;IC8(=^FH\91c6;+->^3D\>\-@UL;AKbc9(+5
CZ1-AI4K5E]M^1M7Sgf^1LWQ:Wg_V+OHO\9;>V6g/LC0QE5YbGb/N3:9[4fB,-g/
<>a[gfV0X154=8>8Ib.W#<S^EB6-^I4F+Z,ZHOH#J&QaKT^V,&Z522RCbL+0.;3g
)Y#_3@VI2CCMd<B[;_ecP4=)M2:9:8(<9OQE;I.7]<Ee[-d?115cK[(LH(-_@HC;
2Q\>a00-@F#;)..5BeeQ[OT3>10KL:<1aSMWKB=11IbQBPFfP.aAY&:X-3Ldf,:3
e:gOA8ZKQ;[aZ2B+7MX&_])2/D<2GR[J)9:+L-]_26AI:/\A&\.b[(/N)T;.^cS/
IT#g[7J[61;a2;Rd-1=Q^J<0dF06)D2KZPP(d++fTX_TM\Kd)SH;19\97>S,>1>W
@DKP8:NS5SCQF6530/b\fI>ccJT^E^22U.>C++3<Z6DE=(F.YTX8ICQT)D\e=acT
W?I,(+AbR.0:[\MeYT7_IT/)8:dUF>+XS>#N)W4^NVU@dQ=LX[]1DNI_NC:,)JM6
8K(GQ@Y?OC9&>;K3Y(W643gPS/&T6=fIIW]8Te^.WF_A?3)dR?EX[0fB@^\Wed-9
Yg:7Q#^^H?[Bf[4^9-=Wf^a00gK<D,7XA7&O7Vb]C?@Q2\E+LI]\aQH;aY&6BL9I
0]O5JZ5JRFUV8bA;C=.E@R:33S_g1NdP/C:^a&5REN1D@[a@--9CV7Eb^I2-2A1Y
Y/36+/A+\8?[g[0O=Z=9J:JP:eKR4bXG::-L<8N@FHN,;M[L@=I(MKTL?)-)IV=L
f[M4=K+6:#R9\KOS])@;OVRdT\Z:#D^fFG6?=^DL,[OE50?YA&=.3(:De(6DUM0^
DLY.dfC;LOA8Q6_+H)[LDBH6>>P#FR8X:S^N39&-HV):694FZeb]NDEO>(9aWX>+
GF6;gA]=RKL29UUWG^Q5YI1?FG/\ZLP+61Y(G+E5HPDY[1J\(]R9>TF>^MJNI&:^
=7)Q[/J8W.NPYW^H\22<TE3e4(:JV;&C?:6(La1G)]DK.>B33gH?Z6/6.AdUV4Q^
gY<O+^dRHM]_90b[M2+6?,I^4Va0CHJ&TKD]X6Of;VW<WMH6^T93YFOO686NR8=2
>\(J2J8MMSa#I(=H-fe&C+7b=BV/RO<dDB>HM8C\dI:,/G(<F26QdKJ)fbRfd]-\
\7Z.A28HF[G;1D5DU3\P9-9MY.]g5,ESSD-e@S.[N>:C0Z4eO[6TWe-fHCEGO1WX
)P<Q?0Q-de)EL]132I&M:V3>TSU3X3a/67aa:G594#IA^BAZcY>.f=P[e_/#0)Q4
=[[(R)/GMD.5,2^7#Fe-)]V^<S@M3X0cX6+Cd+Q57S>aH<6]HCN@&Y#G5Md0fXb5
S2K.gC7N9=,aK/PR2Y)Qe1L/d-[bcXF]//=;5FC93V//+Z)B;V__,,4OC1Q;TbX2
V5@>cV5O2TOd_c8^&IP(O:3Q(@aMQ/-IU;_MZbJ=g5\,:A6&_Y1AaU7KVbdeR-VI
[0dOMA#?d4S;Y=7_c39;)\fXc0KB:ZHI,PZWV_^4aA/MJ7UX5dQgAD82&0N+==2_
#;B;OGH=J:/DFEc=(>>d7I]#T^@=4:&1/-FLeQ,gNNB006d/N/KIFESMN9E_>HTO
MNeY/fG31:+YH05fMA_U3/=OY>J)A.SAW,?Y5)<8GR:4^=WLI1S1e]Ed(e_@O#a]
(=I&Fa,F&G(&;?NA(GRV&a>[AR+09c]EM7bY.(WI?HQ<4VbZ2S2QW.XQeN+8,2/D
9B6;DK8HB,<Yc=4EdANJC,b<?1#=MUH(:GDG]d,+dL:=Eb+-BR,2U(=NZXg>AU,/
cSMWO>V].b0-G-DBIBCLW1g_9M.fBITGH9N0OdTC53:1SB&E,c7@Y_D50e\:K9(5
HfZ,:UAB>65W_43CJ^W?TL<V]9@?@Qe1-L4:X<D]MS0<2VHEBN1R563IB6C?(.4.
27G_(XG[0^HKF-RTTC+G+c]OgR13M46N.O]?/7D^;LZ>V)DFIT2Ab2WcXe]gg,d;
QH^Q]@#[C39G^S5M\/4475J45(BI6USQg?T44F[S?Q,A?FZ)T@Fg?4:0(dIS[Sa(
71MI;=3G/XJV&>a+JdU.bf)K&B0:@D>f)?_ZDCM7MT&(]J?A=D0CO7UZP9EcLYP\
;/[8]?7(EgZDIGM&+TV?-,:KK)fV#OaRY5ES@62P=;ec45JfFeVe:9:8X[RBY5WP
#Jfb^^@I,INc.RUT:<g.@H/+fNSZAfX77L-2U5WYcJUEcL;K9=S&SW(IV^>5_MNC
[L6E3TD;0\DF49;FRE]H&KPHMRfHS_^f0FWT7eQYbX\dK^R1NXHR+5JD^75>86?-
X+(db8BQHg-A.)FUM?<NXE=3T[91SD6)DGfCM+\Jb,<e#3b8Pc\d]KL]O.b6b_/3
QBOT5C9.S9[fXDSB8EBIH[88IM0#9@5#c9/:29(+f/KdJ>dBU?@QM^ICGOaFG8X9
HcCQCRF).#/BU4aTN.]^WP-/ALV;Zg6F0F:ad<>)A48/4@5#^DG\KB_#cC@4OR<H
.CBbJYY+/Y4C1?X^FNO9<IfM3G9O_Og4a#SfP\0Oa=ODfUAE7E<+P/GZY8A2;eEU
#/UNdTMce7YEa3U\WSORJG@7I4#MB5^O5HOJ:e&T8/)]N+;d[5@(dSOC0T<J-LXF
-I=68CIN6]gT_L^_3ac=C,TV\e/^VB5NI<cN5LXLb;MJ^NH7gTd?\,SL/9[V_H7b
F98TJ6K,KJ:UT@OY/eI_4Z,(R.51HYJ;_PXFcdGA.gT+&;M@P8]_V;KMW+U.CLN.
AIYOB;a37g&ZSgJF3A1^O.I5TVEMK5T3+3QU&>3.53OK3<U]g8L^/3I7U2;(N=Mg
VbdK-GT#\)g.5e2WNLHVP?B8,-8]B)B&;_c6@G;G\C7_/KgR39XY-YdcF][:.R+]
\1HN&:[NC)1T)8GEM5>]_cN<^W&L&>V;eP3OdHcP?WTXNIdK1d@P(6PYE(Fg?Q)/
8(O(;a<,<@OMXLMO(@\,(_g?Sd8ab?W6X.eC\39/ZDE:A=R:_^G=O#B/d6AT/Q3(
9<51NH3AN>Y717?0]d.0RUM(V>SU,>e.U-OS_7@8KaC#bP.g=3gd4H7(RQ\^1U&Z
fL>,VN<ee(&@=FD-\bb-P/B/>9WRX6IZ,@WP,H<75GAUE7a:I:>SUU:F6b.>SP>\
-HN0J@6f?4a5IZ/IF2T>=0UUPfB^EOgF.PI]/J5RAD._#F3QGD0e+4+IB>(=BQ6Q
1c&TMVeTW,4c=[b^PPIP+=VT<T>/YEcO6XQR:0.^PQ0>,=L\C#]bN&V#-G.-cRMK
,Q]8ST7&81(#^0Cg7NQfV:<W=T2Cf;#9&XXAA7bg0TN7@NeAW/9_:U^B:NT&a;9D
D/3aQ@7XXOP=QGf_a7Ke=Lg-WKNX_H7.YcCFYA6&gH\IJScgL]g66:#B?O(HWU_Z
QC_1:#7^^R#U0ZXD6=XG9(FV4J-)9H1H?TD3eN.fFEAb8K(ZQO9EgS9#JdL?]J-^
.PN(#>4AT^I.]X,N@IUc#O/4.ZX-5cZ3AU0)G9;fSNFDZSf>AL\,.]]V&J5GID1e
#6&0)[A=<;JdF;FN]]@?Q3;NU(1HVKE/&?KF/:fcgBPI)M[:C#0C1DcKdK.6V-dR
7Jc1VV?M8BZ=&\_6]TVa1)^a]08@YP3fL6/8L33c:Qb&5X&_8F=K=IB[3K7e_NQf
F.J7A<E^F:I:cb^dMe]A;C;HZ5]5CCR]>:VN0a_[OSE;+3@aWTMRb:#Z;+]P7c(I
SV&KV;&2XY^[2UP[2+&[CeBP.L5(515MFP4\,V=:;f67__&=8_d,BW9OFTJf@SO)
K27\QDAGD0e8#P#ZX9\eO@==&TMfe[&PZX_N92b]PZ2@eTG36TQX+,IFTL;b(\MC
30C8J_T,+8)I^GMZWRe740,0VUZV??T#\a@E8#(8>7WZgL^L-@(20a(#O/GFK8)N
3fZfO?ZKN(?Y]=>3&P[E+[.V;T\;S=F1(=e5bU5F6MGCDG86A19AE5U;K?URSJ2B
ePREK@eZ;H)/D)Z=@H4S0c8_9]<JbKJI4&&GJ9/_6/#8#SHQf][TWbL@eOP:IV85
)QSE97//^VE4Z>=ZM<:6&/-Vf=H@P\.EUI&G81@A6F:+TVSGCI/^18.ReAM).CG-
Ca@MC)YU:8_K@g\F<5Ig7#/\b;PJ?OQR]YM[BT7]JNS\_K#A<fF9VO=b#7DR8bL7
_CW7XDc-dX]@KEUBCRR?ACU-fMZKA..H[4JYGKEfNPMb5eX6c4a.==aM@NR]RVG?
EM4(Z,9(;fQ.R9AMgJ);]F#U-=gY81_T0@_RK:PWA,FFCVgXdZ/1NBAVT+Y@cIDe
-5Sa3b2:<Pd)gWd[WU;]b30J_&K>GKdI&&@gBU7gNJ=D,,B,=_.gH-B7[<EO,36<
:Z-:P@YG5Y[#W^a2B,HJ?d-^=Dd417gO-Y.Q9PWXX=^GA>T,<R12cG>@CID/a<>8
3O78:?V[gbcJ9a^.e1+MV-7^>8b]X>9YbHSN#JEQBJV0CSVQc5=/6Z4a9ReVS>Eg
V<UAf14.MCTD-Z9)e=_PZ&PcPa5A2I_O],TWQPWC1_LUNXQN^/UHbQA+5a]J@E\C
IINW:5;+ATW7Y>H26=;]:BJ.?aH1F3B65b]c@BCV1ZG#&J^6c\VUW=J1)\a5QEXF
E.Q&<].8-@+#a6]R[OB?MA&MFJ)7J0=T@MM[^b>#^<ba,U<40N(P]f&NV)TU#gTg
g:([8e8Jb?5>\SN,Ld50Id/<(Y2^a,6b@&1?=AXOOFGcC9SY?]H8T;?FY-?=VMB@
gJTSPD,QTdBK5>df-8>0>@gT-Q@b&gG.>^>da#IJ+UOA6gJf5BP^OD16H0JSY7)=
J(d=L=W.HLeKQ\W^3\ZSK2@O5-&gMcTb1ACIJE]I0D/DBW@LDJPP-;??:3U681:5
)PBP?F2@6+V<27cV,(@><P(DR)QU=IM_4JL1@NV2]FgE@]_KR63DgB=KcWF)>1f+
S#\KF-:5,&#/\M.8+9]>V&Fc+3V6NFW+:CUYbFf-X@GYI4WKG]P1Vd2f9gMA@B6N
1I7#WcF;eO#_V>1VP]1EXcLPRMIU506\aZ@)XL)<0;;,YRORC[TUX^J)0CBbOcJ0
,97<CKZO([39U4F\S&SPUeT(26fS4+,@WC7J21)B#M^UB\;Q8^_0/;EZgUQRQ<HQ
6=U]IAfO841Z#^V7NCJO6Q].4>>SUJ&1P@;)]&_HKbHXdE:;aOcY]3?@gKQFV4Ib
bZL+V8e)Zc_W=a^eV7C)H&>KGQC@^YGN(2GBN.+_cfL0APN,CD]^Zd\gSe/U<R>=
ELK;;H&e4T,FGe>:4FWcc:]E=EVaX_VWG(?A[2B5D3T-@61]?c^[9Y=EAATI?D5H
.FaHS(,DF9),X92eV[-ZGD,1,VOOVK,CEP1DEfKa4Ha;LGWI/9#.b,V.><H;TG^D
b(W.XAN.f,J<Z)#_=d/_Q_XeULZL)/>IRD0e9V=-ZC0=UM)M72FPeM8#JC,Z=SEH
,e5W7VMMF^=Z_e5L?417[_59f3&1F\>WcF<5O-KKO\T@Q@[;^#.1-D.^b15VTSfe
3X7ODe\==/8739;cN0Y3=:ODdH8aT8/2JK?G9WYF+(Mg?4,=:9XR=8+T<c<7J(0A
_<J>DYNKd;1(f&S+(^9Y]=dLR/DZ9519fcWXEKCZR2YVN,cIc:Ld):,6A?4DKB08
D-f(P?EJK+CbA&,V2c6N[6.\VeFgNRFS3P3ba5HcId07MVF=+NY>N;<,LA,8g@Zb
ARL1<T5CPH>GR^TNb,6HSSJE(RGd&?[ANSQ8E[SXXS5>P=74g9IN1^R+(=:560BQ
TSZgT)VOC;B^DST[:U3bPVY+ML-R9Cd/Z/#[@bUH#EJE@&P-b4VMW<4KZ(TT1BMY
c6LDQZ;D6);Dd:Tgf#42&J_J7Vc.9C:F1GPMc?T#MY+cLT1H1O82]Fed+1ZD.R:d
5a6Bg8N?R4Q(d-eXI8R3NSW;V/FF[\@a--bd6#b?TP_OWP4f>+8?6W/aBSWUWNNQ
&.+eHf[HbOW;YDfL@--.5G^fbLS\:UM)fb;R=19Fe_7TP2FQ/,MY#HGQ/.CBa]Ve
?1Z1B(&J7SCg+c0.Y[a4dSCJ.9OS3C.F@5Pa,+E\@UQaUFMMbAJ)DF])f(H]1Id&
@(7&ZeG0Z;g@efY>2cQ&@\QgeDbbK8FdTW#9?_B+&:M]-M19eVJL.-YAV55(R-XP
GGS>T@^aZ>,B&gW;L8Z7V&5GVc0aV.6K01fJ>c3XC_B/eM4[C2H-+@P?OLG3I#W+
+A)4@?&NO1gb<?8g.]6CY(>]0NcZ9+:(6?H-1&29@^)6G^UCf\?Z.)C92/Hg^ID[
/P:F7VO0Vbbfbb.Ed4dGBaV-gM\&[/89cJE6#)H+<3^cddW\Z9@<8aKZ1897X5(X
1G@.@34Q2R?RJFbUa#cD6K]>GOg^<Z\>Rb0Kf>@.U6,X4W=C?YZHD4-OV-[,/#]1
<RPc#N;LHe.V]GGMW]BYSY[G2([PWIU=AfW=2^0Tc1&8Nb4LS)_(g_9a^JF[@Ec5
?_/fS&YQ;O^gcGA6SXUXg_VddXD01,;\b)U4[.b6]d7:g?Z(cf10-43BYO1S\9>8
cUAY)J;?LTf.TLZD,HcT.IDXQ??882R7QC]3Y6J2<BbE)2UXW7ZWeTBGSVDA-6@#
QS?KVM[DDG-Fb9BH-F)Q<ZMRF2\O/2\JF;9Cc#^M=f#MZOJ\8U&5bOT-@E6Ae4V2
gf]:>M/f99GO3MUTT=HAe,8V7H)Q>\V(^.8H5f-@G&R>GC,39O_&=79E8fB/Y<Va
9\\@5>AdSRd\A:@J6_IcZ_OTE,Ob2K@-T6A[CKgE91fHB:b(d;N6Ad][F:?^8[6G
+B6G@&f/P<LM,#VccE;BNW1^4,/8<H3+B^#aACW#E7,Z-<D+/+6;P>fbQT=H4Qf-
35(599f1?,&Y8X?<aZg-e/138UJ(<WMVQ62J5D,]aBE.&65(??(Ga?UW1T(92+:P
;I+NH_M9f:IaAI[gc#YKL9781DZGc&R.^McULOVg;21AKWaZ;7I:-PYOY/21A_#)
?5:/fB#dAZ_9/-&RAf=RAB=P;64S3:H#OB:d0]4X6f_1gD9>4);A1]8dd^1Y\&;D
1;Xf3gV#DfEcB0]&.&BC(Q?ceYQ_92X2_Q0_c>S-aXAW\f9Wa\EC.g_ALdWL?;+;
)3<)5L/Y75#&^>A14gTP5V.\e+^EC\&W+Z;5#6CY&:58(+aLK<AI0=_Ve24<8X<+
FMg1>dUKZ0bXeZgg@e:^L&.]\7T)O),B2EWX[9HCaFC-Qf08&49Ud:8<Z.U8X2<@
EP9.<XN^#-@G&SWJXK+E:dGY7J]^b8aJ95&7a\+eDdCJ>:f5W#R(,cgI@17L;&?G
.:ec6RM=Rcc9EN=I>_EaJ--8@,Ue5.]4-#[T^@@\O=JWNeQ+?;9_Xe-EFYD>fP:S
DCZ(,b5aS+=MR0A#8gJ1/X:TeB-EMK&-e:MG]DL=7;D[I(=:>9Zc47M(35+6[1+E
02Bb^YL]A(P8L7-=#N=O82YRU)6CH@.([MgQXV=&2;/(MbIOT]6D@cDA3bCE&0M2
X:Ya+gQ<>U1<W.Ve9:#NPINc-)/.70,46#PFY3H@@(@Ff=SK)F<?/]]]f;3))4/@
684@Q#WB,&M8.:CG49S^-G1:c4^9[@@7M^EG+gd+]TdeU?X^DO])BA();&gQSEO;
-BYRRBU=R;3SI?(X@&0)d?<JITUYb&20Q_-2<\GAG,1+0REOUKNFF:0&O&&UN1Ne
MQ\_.2>aN>X(2CfO@;VT?d<APQ5:V>8F3F6S^>#<Y\[#G^,-P\dF1\\bAZ&CIW8@
e3NYKgFHJ2f;&CcY6/6KPQ3Q1==P,/^2b4.0c,UXd40=(.64-O\+a(A?_@/+X;aO
NYeFWd7_-(DGQOS5F0(gPT2;)14f.WMJYQ#>cJ&@\e4C->X>J)dRJ13653XeAKJ4
e4C/)bWXSR,+6+AgaM<?=H4V6F4;a]a&N)Ng(O5PYTKb8AQF6YNXZ0AXNb&O8&eB
NIF==&CU6e>E-NZ4Ud4bT(0DXVOGc1UC8GG@])#<]NGO0WK8QJ24a9IcO_I1]8Ma
X;aB^4)fL5J_e0WU[bYY]#d.gNHD(4CC,?@<SQa7G]L[Oa7IPT=8:,gDf(>/V3Y:
]CH2LC-40=-)M^GNdS.,Zb6LC\gOf.NERU;bAEV8g0BXX8;8Dd\FMTTT42ML[C.B
7aJe;WSJD<:?\A#KTC].M^gPGO6Q_//Q#c6+M3M);26ST27ZGGM&(4LU)bN>>cFM
>([?Z\>+EJD&<WKE?acO5P)O7AC0=bDC7(-(H\XN,S08U0PaYN8bVA?U+@_C-6Z4
X4DaXC<?GBI4=VV07VHd?,81FB29?]CF=N96?(&WU\F)F7GY(.?\-S685G@^UI_P
2WNK5O3^?)&M^(#L:_?4YF0?]#/<V>4AOO#(^FU,LY/gfY&HJMIJTc;FQR+6_S_O
&NLHb>+W?I26GFES->I(O>VJS1(=>WL.=NTOg8YYY08G_N3^_0Ub13D&eG+DN0cJ
/@Wg:?cD#^XJ_K>]_1L+QWV)?CZT:<g@-W.&OL63P):G-dB#dBMgFbX_J6AX[DOH
)D?c<W3M8&ZJKcE)_Og0g0MZKAT9,aED_W^6L/.KUA,b^bX25gS]WMgNW,\O^SHb
07E\?LP)H4R\39Sg8LK4ZRA-89GN&()Z:301R[f4>A8-SB4_Mc(<G)GaBFG-:W,5
?874W]PeQP0bJ)SQ/+52U;H3H^>9-OdTU>:cZJ]g[b5?a,(bcaMYV.Y7_[?8/L:&
P^e8=aI[2POIaG<QI[ebO)0M\^N1BO6:-JSPf)IE@e-Ef+-]I79K\7G7AIJG8QbB
6-B_OK,J:V)Q-RW61[.+Ab&AZFaS_e+KK=5DBG[bCMA<)M^-cU14T@(#+TXAe+?7
>W5?W=;/O\X812UVTL1C:P,O;\5M:B?HVZ]N^-b:=&[_]_2QT18eeAPGBDC<IS=E
Y8/^geg1@e@5OX2[5If(@PA41VDa8Q-QZEG9RJ.-[HL)PYR^(&&(+H(^AO2N79PG
Z>OW[VQU39(M6&;?RV0QE+5fNBDgG674G=OV5c6>S2L\b]:@ML&=aB,&[R:J045]
U(7]#59a6/>D3g3dO5.RGX7,M&F61F,SW6bP0K(V@XgA<a6?L>WB:7a2[AJ+(92V
N:)gSN9J@#JK#Uc<H,2B->V>ZCPAEeRH@;9I7eNAU>#)bLG1H6cD=.E[2>2=2)5S
K33@+X9R\K7,B9f?^XV;Ra:<T@&-U]7@#UPCg=G:V?NM;;(3ZUgT+8BfE+UP<258
cUD?S5#1W=H5QHZGfB4:JBbGL<IDXP<Xe6#7&->99:C[?8C9?eQT6+SdFP^JLX5-
&FHG6RZ#M06)Z9EMLAd@dQJMZP215F1a+#&0:0L>Tc8IDW(Tf52E[_LSc.^=D9+(
?:Rf69<95aC]RV^:0VWB7G=N6BbIYDNLR1YC#/9CI,/8.DSU;J]..dLOH+gQAQ#)
/TOCGU472I&IV)6\9\-B,;MHdUX^-3gdET0RJ4C_]H.(M@<M=DX-E=Z&6:C_^=(.
&.?3WY_X#d+K2Y;c+)U\]DEB@CXZTWWGf.#=H_1Y\/MQ(0ULe,QY6DPKN<TK1^MP
AQ^g0gBb?ZPF8(dNRT=G7eH+-A=<N96FA[6ATO<Sa:[+Pf=I;<^V\B4?Z482f.#D
4J7(?M3;OBT[3,WL7QEO5-73#EE2+YZ,I;#W2O79f-W2-6(OTQ6[H5,B>6X#&IU2
gR/<bEgHQM.4^cb1NDa/R:FG1c?[=(:D&f)?(cX7X[0,Xb1?YZ@@8:D95<5QWg,-
YDLVU@#J;?3?B8gMW73.;BbX(f1P=JGXJLG^NS5(K_/XJ,6?aHb6O<3X,cIAUOL+
]AfDUX6@E0L9KGC<e_FSF3OMTBbDBN[KGA=2KS@O4Z#<9Be8d/ZF3BgBeaA0])[\
4H=BF>c4&e-@[]>UN<#>V3)OMEG+-15GB^E=CfA;fG.e&ID8)E;gEF(YS<1)a6>-
=L@0S]bZ[H5H:W:bY[.8C/;D\RJ^=^5TJ;@B<-\66\Wb,GMf,W/>+P^8(PNI3UZP
R&K184SE-_9-Q-EAL=HPe&@I=(8MXQe:]OacB_>21#Zb^U\8+J=JT8@D?U.H&J3-
XJ;LDZ_[[ZP(S_U^O+^LGQ?=RAQeYg,/Z+0(IC+OAXED9F8QAbP-^UQag2VPB<63
M<Y20L>7_Z[T#ZfB@_+3^4P@@Cb+DBe,;:NNHbgR+GM2R@FN,Q;<=]Pd^J?<?GCR
F+LBCa8P8b,fZ8C1J_d(J+RKZ[5c;&G@G3XaZ>+XJfF,6UVfDHXYW(?X=.2CG)5>
KT29H@+QF.4&F\\EKLB?LG02IXP6.H:[Z33:#_>Q?GDVYGfd@AW=\S]@.;=.]Q-c
b(R?fg=(B^>2GCGU2=(QSB)DZB#-_;PS,AC&[@&G_K0>,Z#)6AgB:K3M^]gDVc,S
C^#//,=11[V[_Yg-^>NLa^9AP83#)R[Uc1,_6e3,@E\Y+Qab(d3L6CLM)WGU<)2g
49gFg_;\FRDX\(SVVBQeg^gP1gY>1#Y/D-6G])]7F,/E&P1\dd-(1RcY^VQ(&6_H
FW?G39CR=?4P[7G4[E,)Q-Q6ZAPXDa4@I(8(RA9a.Y)2#C=VY>TX/<dEPK+]G[KI
J@#G]7;1g@^<:?\-_LDC3HY7SDY_LG+X,@g[ec>-[J/@W1U[M:-fDF2(0./JERRH
(N,:fRW92.48IZ@8<53XDa22++OL685W_WK#b@86PbTOg6F#<7ICRQ2Z-SXX_DNI
_7J9JE25Z:5R6W1UZbKWQ<\bI8W&d<]WdWOJ_fcN7;(E=]dca,&0)R]\^dgY/geG
3dJOa5cF=d[ffUKGMgb<V(UeG_:BO4V0@6B7_(ed(1eRCY+f=7+TV]&LHfc15JF7
4E9b7c]<,>Z^ZeY\4AWaA4fCZ]g#@T\@a:g_3N;>)2T3TN.:M1>e4)>G],D3Q;#+
Yc7Z?W;bdSI#.#0&MZ&BJ2^,5Nge5SY/fEM[R2W_PfF>[2NU;R:7]RJdbc_QEKUK
#>@_S+_#GH8JL+YB/6AQ-;eFe9U_[\6[;YWN,<7<4DRF=HP.aWE03LcEgGcHXJ1D
a\=d>ef<5^3S)+9GYXHb][8IIWS6:aTP>54NFPNJA1:A.//ZZ\UD.1UVTC[cKZM6
XXP,Le;KG^NCJ=T-86cW;H>#[V7(VUI[fZMCRADQg9gRQ\E0M,&GT5PDg)I;ggSQ
Vg]==][GMKO,@f\)Y#7K(_@B0.]N6LJO3\(]3.EZ&N(7S-6_T^@cU>PXS]3#\eV8
:gcW(M;L-DA,cL/#.PfVQb^V?Z024P;=ReF>NWeR3b0f]?7g/M]>ad]Ga+O8?R1Z
&T^W?SR#@f<IB66O\YFKF+]_92-37FHM24T>1Y?^WJI(:.DV\QKAKCL=gb/]-E]f
D[K7g_,H(OKQ>P(-=4@P<V+d=\<cHQ,B0&H/TVZB@LW_>Q[;bIe,DYG3WZB69@Qd
9&+R><Y(YacSO#IIX<+?N@YU3.AU^IWJ_Oa?5D@W,cV;CN-M)b3M@P[XWNCB06Z?
^f_-Ke/4?K5)(>&DgQHEYSA<WP?dX[C)bMD)RAT+,+dJX0KEX5A&YZf-Q1DMgA0F
LgGQ?P)aGXZ+=NRTYV=Ab(0753<DN:&B+B4W;LBT#Y=+8>#_+GNIC-B#5UZf?[SZ
(:@R0789L1,^1NRDJA?-8FIG)BPR\Ce<WABU@9C0AVGK,E@C]Uf84=[MAcg\N,:e
6;XAb,dgDf=Ze)?Y9RSU842;#/Wg,@\H;^HD]2^Xe0Ab8_563IT((DSd(7585U])
[NR1,W,X8NBN-L9PR:D&If+7-E<C_@IDRIZDK<PPW&&C>#f=Z/ORI\5c(=UZ),@I
I2?@E@W1bK?aA7:QA-S&O=D,Z#B0(=c01E7gR>0>dfHQ(E;--DXFeYRYUCP<KR[8
3_3N3GW<FNF:067NGf<fDP65ZMQW;Rb?H.PL@U)AL(&2,GJ7IV4g2OYPXV?E5@=#
AT=K=&S#\IF^c+dR@HaQWYLJ?@J,\6@0,K25?M^Tg=c9.48[:HJe\RaTVLW(;THI
T3YbKL]417@-24L8#G&:1S,]?0_f<fM5ZJ5f[;AKL5(<0=M-R8c9fRYI9=e>&)25
J]\(YQA+J&P&Ub#84>TaG<P=P9ZRS^:M4LIS)I2[<4J=a:C0M2V[FHV</a;c1\>+
R[V<Hafb=Va=QJ@aT=RKfCY39)?,gc^Cg#EI^O@b:aW]Pcf\#I;:_>J.3\+[=]M)
c9TT1&,AFLJ?^\]ITS[FDGP]FgAV\X6I(>Be;]f6KL(OTDEd-eQRfPXf^^-2@83c
F3[HBR7&C=^=]d:HaTT)f;9&3VNMG6>@He[>#->UVHPNB7\/)1]#JSYKLaLATOP:
@(<Y1):M[52fcGXJEG=G/Bf449A]TaA(CR2@;_]^QSV87,Y<(BJ<M]P+eaDAQVMV
#W@QJ?&72RaYR1[5)5;aD]O\7g210^7^\dNVFAQFH@Y&1c9BX]]g]]b>M9V:D(.e
ZH1f<K]+VcQ]:f1(4#49ZUL)Y3(+eK4+-^FX@Q[9\R&eK#]F6_84B\N0/0A(:ce:
NP7NC6BOT?DC;ebTS2)S)N0bQGZegXMa6K>XAE0dQfO)N(LS,FJ+dH&43>0cAC5Q
,gUS_gNQVQP=V1H_A@9E@/#Nd,NZ7-\LE,69Nd]^eZ,0-c-2Ba3W4Y<;8PFK6C-c
D=6a-ZIUFZ#,L4LQEbG:9dXa2&MK@<+g1?>,&g=?BRfZgEOfK;QI7dUWPV\1+3V4
B:bF9J72)+W@G9BAbC&5W/0M7,X7cH1eLYP2+I#ILKPJaA8K\E<=LA<)/I5D5?.<
>1);MgCPWU^QF2I73Y-6@Y7X0?X=UJ_.)4:EYdMB;O:Y^[-M0gcEfOE3>N0-S>-0
ZT1[C+Z.)[D?]@;d8NS6/(G+XbeNb^S:#QOObQ>6E:b+fZN,[I[fYE@QMTc#G9@D
gc1gf0dQ5<+PSd[.gNdAaH).E)c&YGc7T30C73@\WBe/E?aRKH.JP[/><I2_dWCW
/JUSU=O)5+Z(B9UH\Lg^G/4+cFU2D_J4SQXCW+Z/Fb#[=TKC[JBM=(3g]3\+]>Z<
\_&<f:715];);b5Be/,E-Z4(@:ZWO^S+7eV;g]MI+>VXQ0?I-J_TGcc[)I9dE)KT
CZD#1eT&QA:LNKB-=2].Q/+_aI,<Re^I&edd##67XCDcTAHcQ[6#PNEfC_aI(AJ9
N8DS?TBPFR5W5e&LN8@B8J>>T(\RKMa)BW#;/O\K8A4G=2Ygc50C:(aK]K#8^_5?
#Z3;&S5:[HLFa,ac=U,HVJcH23(N,&I^0\Z<.+-,,-D/3E(//=56:HXJ0HI98;RO
Zd0/VLJ32A+YJ>?V5;>-:9IgI:Q=c-YCM9C/e@F]/A+#_@]BP)R82cPMT:aX>]8^
NM7L-P9b^I:@(OK2.@2I)/VG&75PXf\3-Zd)95,df==;R,SAF=-OfG-R,6R6a9KR
N<d<6S3D##Kc7be?YCT59V@8X>QXO3FOY&YSMeQdXO(D8a9?[Lb?K93RbESY)=,D
A(U#0=3PYF#CT\C30gFDVPX311P]AQRUd?Eg4T31+dKDa@&f#7aELE46f&X;AC?1
@O?[QQ(=U59P;L_GOGFc[KSO4T<D_^.T2UUI7/V9@+4?RA,U,+07D<PgV:fc(=-6
L#SL2YM0]fH0LEVeNd[]5S?T59H33Wa4=7_Yg<,&Y.U@#N=E^>]b:g33&)W[G;L<
O,6^#:ZS]B3aLJ@2Fb[?>_d(G?Df;U6P,6.?#I55NCLO((M)F:#UQ0IU##0gV-6[
_W;J;F)RVX:[KK(\&FDB)OD+(RG\)fQ<ddB^=#aXg]d>,:H-e2SK(K=]N,XQXAAK
]<MU)3J0C75Y>0A3)V+54\FS3_8[R3a7L=3U<8;?/8X/G0,>/BU2BOQ+a:)bBGdA
+<<PO3DB9/=])8d5TTAebN^Ngg&8gOU^;&<I>\JbIU3V21-^??=8KHG5JW@B+D.N
G6dF6O8U4;gA.^W_Se44DL&;F8&/JBSCO@:BXE,NdP-JBRPc^8ReK]G([&D-AL?G
]V>))QEEDP5>_1f#f\UbC&P&IYWJ;Z.,>]W9?]A6V3.,>&_e@;7WV<f42YK6MVAM
dPLOM16-c);>d+-dG7OfaP5f:?SK8>RDLg1=O;H#V[ZG_&+-B;S=D4+T_FFVU#S:
_WgF4W4J+\9>9QLM?_Y5B]_)>Og?++A?)WSdN.fQV8g9.T6NB=8)4[YJFKbbG4eP
>T4HQR0ET0>+U(09/<=Gfe8a4<JDB/WfH8fLIVPGF8A3>C[I98\89N@fMaD/N&E)
7=0W;0W>ITa[ZL,2U+Rb/DMFY#De3E?\6EYb4SJ>HYL8[e32HP,ZO+TQK&M1IS=;
C(fA;_>P+\aN>UO^^+a:eGT[X/5>L[e1WM+F2ML,6V4RS>1=)8V-2RML8K9UceKX
c?:J[CW.:IYQ&<5]Ke#1@4:[QS+(KIRJ)YMN2(RbW^c&+L:[3CDFA3&S5O?@/R];
FXgR4,<FMca?4KKN]E2&KETMMJ]f5Y#fd.;QTfaMV)^Ig53)RWCW=//@BfLGJ5-B
RbKeTXYMdN2+YdZFf@8SY]-,KMPbNR;[E-.],&_R5eUf=+T8;>\Z#8A#>&1-D>\d
X1XS5=X8Q]R+D=4_@gI\d&Q&-Z-f@C9JN_E(I+EQJ=5b3McCKdDDCGbgP:gG+7TK
cP^bf7)1GD?_dJ)c<@NJV-8)-80JU=GW1ZVc6J6^.U.bL@<IQ8O0.^)eQ-[=F.gW
@?D<IX@APZ11AY;ML_FaScaTc^T4PL^,L8gKdf(KIJQJ+Ef6d-].?DQSgXKPfcVD
+QdI,[A/R<MVgW3_#5(MKZ+Lb8KcN1SG&&NRZ#]HRYS2g1C)&g&9YSg@3_SAE_?Q
0OC-,KSNJ3Ze71&NNd1)aU(&KFAF9IW9YfTHK+a>G[f-(V,,XP_LAL,CPY+]4([3
YF7b\Y_RX?H#Z70W,B_#]dPPD=WO?&9bR&d8ddQ:7-3/&cBX)+WbfbfZ#D)T2>,&
<L?3/A(ZZ/cK/-#Y/4EB,ET/67#)M;2^B][,(H)gKbbO_(Fe4[-&YfRa];UfbCOW
FZ>25b4V^GDB3a>>&f:J.#S3&6J=W4590-OF:C4a5W=14,1JJHW.YV46;cfGYMRK
eFP);Ee?eeEL:>G]fIdB.;[Bd;F?02/^\B+;2X@ZBN#/[b1?<GBVP4:E_F?LZ5Fb
0O-0RGd?M:2)ILebIdcb3=V]E;JEg\7PTaG8M4O+dCeO#a2<:HKWaKP/b2(B[Q/I
Z#@EQJF0\5cd4C<@04a+N^4JYULC00+P0G-0ZYfY.[<M4(La?Q^4UNC=V^F_R2IX
bWH6R4S914(0S:D&LIJ?2D&BK23&O0@cG>/?@)</?#K?U+aZ&/_baae)TaKd>PXa
ULN@dB@X&[.g^-T9I8^TE6?1<a@ELL4g.UgM^#:K29[N=#561gO6\KDbCL\12ASa
Y3PN&IHA^I/]5IQc,dL[P1&)W/J&WKEPHf=:A0Eb/Tf21G:/0\?=Db8]+TP26)c(
c]_S3>NW&B93)3H9K2cOIW\+5g8GK<T@K&bc/TE(f>&KD/a:f?Wc<_Yb#;1_AUEa
<]#NQU0C,=B]><eC)=ZB1I6,]=ODY0RfdGTK/A-,FVTKH$
`endprotected
endmodule

