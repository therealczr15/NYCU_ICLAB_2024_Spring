/**************************************************************************/
// Copyright (c) 2023, OASIS Lab
// MODULE: PATTERN
// FILE NAME: PATTERN.v
// VERSRION: 1.0
// DATE: Mar 31, 2023
// AUTHOR: Kuan-Wei Chen, NYCU IEE
// CODE TYPE: RTL or Behavioral Level (Verilog)
// DESCRIPTION: 2023 Spring IC Lab / Exersise Lab08 / SNN
// MODIFICATION HISTORY:
// Date                 Description
// 04/06                SNN Pattern w/o CG
/**************************************************************************/
`define CYCLE_TIME   15
`ifdef RTL
	`define PAT_NUM   5000
`elsif GATE
	`define PAT_NUM   100
`endif

`define MAX_CYCLE  1000
`define SEED       2024
`define DEBUG         0

module PATTERN
`protected
59^EVTdTSZE_EY&K5@fII657<5c\a=&0.bHPfEN#ZJD@]G(,^6U],)\D&.3ABN@N
SaUC(/aBMI@+)/KC14?<:b.@>-g](a&5.[:#P.:>]2aYa\Y7a7C>;2[;M+(O,L=J
cA<aV7.5^Ma=27V_<bY&dUK1\>H&H;SQ<FP0D(BOKO_Jf3Ve)C+Dcf\D8#cAJV?\
IO7?HY]O1:#gKK5d&)b.NLUE>gLN9O@afI>?/3S48A;fS?EQb\TPFXc/_?5(1IL<
=Ba33_:?g7ea3+O#K6UEBS;3Y:cf/16GEJA=e9?@;/B-Fe8X]^YHgL#_Ef\G0gS/
#ff.3)HQDHTRCGNeUU:849&e#DF9YY.PAH.26<JXFdQaVFD[T-1Mc?d#A4_8&Za>
KQ+^0+a6X9/BFac5gQM]N(4;GCH9PY^SJ\Q@^+[VQdU6JGY91\ZC2S&ALAJ57Z@E
^+L)NUF>L1)bL^;]>dA_7/ROWS+:>.)ZU_4M5d<JO(JP_+&:^e<,)6HUKg<E(O<;
^Pf;Q0250[T.\SAU\a#IOfP>D@J;7\AdNbSfO^;PC4caUKZNL6)aX6\caO:N9-[f
P=3U6=eB.)16Q1,fL1=LB5,fM,JFI/cGa9]SVNBWTVM=Q.K5<8+N-<]CgM=X,X.8
bD,O_+9Tfe@R]O?JGY))&65)X:VW,dFJ=B78(+\3&ODYMJ96JN625S.=VX#F&SbB
#:93.LGPF)RCN_eKC3S;_-)5)Y.b3\\?:eV^T./?^36:)?&MH\P]fKDGJOa2Hb?(
agNbQ\9ZgR4FgC+Je:\S6]RK+6;&FVS#THK5PJ92Z?RZL)7)D=\7O[c/>Q<UU9H)
\?(F73>QU-LF2;VN+CgM7J_&G8=LXSAZW;=8H[\UDD=c&Y9]1>E#QTA=dGKgYCgN
Jcb7.WbTWKTSH>M]@XgIF@+IQ2.:;G)^/]QA6EQ:BJ:OJOdYW5)4N@>2H&+f^b2^
]53-OTL-S00QP9]>);,=K4:;Z6-S3>e1+fgN[_gJD0XBTYY,cB7@(7MSB?QA=c8+
B4Zbb:FZKKK>#\^^J+b-#V+5(1OTQ>21.&Q)_,Y-T5:69[JEI5)A-L,A>=?9[D8f
3XTA62=[-cd&Jg1H?aXN)]dQF?4?+E-XDE44L5d:OBafFNf@\.LV7.ef&CI2OQK]
AgOD6Fa7Q^PZ5&Jf@f;,,BN<:^M:2.Z7Hb&QVA\=07B\:,)93.Y/AKfI+^\P9g8Y
a;.K0Y#_:LEQ&GOTU+8:^S/2HI@M=D3@=B/)Ygg9(^)fA8/;)0V=/(+\8H4b_bA0
e)bI4^-O57IS^(CIMIQ;8DL&LdSXMDDL-b=N0=?QLX70\S\fQ98X08bPeV=U\b56
;&)8MH.2F/(XKQDU2=#RS],/^:U7I@#Kf6D(^AI3_H0Jg4DV\9E+H^GS_^R#]?5[
QTV]1+&1f5S96C0<FLKY.RHS18-aU3,I=bX/f6Z4(KLJI].Q#Rd6KHcg6YdEMM4=
+/4f2(HeW,Mg;VPG^J[,Y8L5@F>[bLC8JT^Z5;O(2H6aPd>E)Jd/43)[M7C,_J67
Q4]g5;EeJ?O92dAbVCI_H/g>>?-UO88U(EK)Ng]79I_A<LD-Q27WN(C]=5<F?#>R
(K]1=@:M<]BGT?8WRN4H=FfK94aTWD<W8\OX.45Hf0./GJWIMT3:(+A.X)b]HJ@^
90I)e;38MXBb^1_L]BFaFaC:8bI)f.I4,DJW<_W4dWd/FR2UZ/C3-e6<>^-#?(=M
TW.F^90a6/NRF&J#?T=<MHJ@dIfH<]gP&d/#CFO;X)BS+K1BUB\MJ@e39Of(Vc;G
1GK9-.[4<?9\:&PWdW90K7=Oa4#?bQS/92B@RTC;@GS.d<+b(]fI.U3B?M\5SU-4
04..Y>.-X_),+[0g/7YAK(3:@]>,[[(fOQX#B/DB7H^7IdUdMV&>;dS,bXH0P_&.
&Ne3#8#>+M@;C@a2.[-Dd:N.EH@X>-6,/_6Ecd75ZfZ4P8fCdV5CUV:gNg<UQO(.
.6@@g/=RK13BSB2V,^9QMNU)J9\dO_YR,CZ/P6c?]QcJ1K^L_HY[dQ2B\B@f,FfK
eK+^KAd=K4Y@CA_?BCI[4b\<_&;<c_6V9SGC,3bcMcC7H?PMagfN9\>LTLISF/UG
b+798V174>MWA(S,KKSea=;#FCDL8SNGZNO^R?_1-><4?12TU40,QBg^^]W)QdSU
2g856,Oe69gLIaFDU(9,87>WP,PF-8&+KXf>]@-Y8;,Qd+[_7^[7&4e^QJH/V,gb
F8P4]3W]e=Z>:LJc0dK^JXbNDEf<@A^>[V/S&)U,=J<@(#Q?=gf[FB/&DWV]Xa)V
UM@fd8W_+PT(=eRJbcd[RC-JGbb3ENXa9@EV,.#(SJIQGaEVTB#5AJN;@=RTLTE<
>f1dfAD;@dcA2eDS7LK)f71.0E#?5R>,IBM3A/4[H4dK@e_0B@6:F--/2[3M-&OO
@UP].\YOW>W0+\;Y@83G#5[ON6Y:K.;6#9,[Pc?dD)5>.;MR)BD==aL=KTcg;;K=
0.[NX-d,P&\T9+ASDG=;N8?[dLLYfZFdCccM8\=EbJ0)VB@.]KWH@@/FEfXNH[JW
+NX?Ce)^J-HK1.1^9+,DVWX?FKMQaK[Mea^;Q_JP=2g/gD8NJT#,#S?V\FUQ^+V(
_)UVYH,Q-^V=0e]9(:S,XM;#RCW6KGO\69OH^bHU\FY=Fc+6>ea,5He=HX;ZO07c
D]>9DIW&eD>_d/K;T.]>IDZcb62@9X2S.G3/--0]aZ]U+=9@/&I3R(:L0E1G33?g
da#7VQ-dV1bgUL8L4WVKF0H0Y7Gg>&,/Tb<A(2YM3BAacdd[XJ@OcF/SD:_:H].1
T.[deW9M\X_2S.1/+O8U&+#T7a,A,JI_(^d8\VeFK481_7\Z3?J-&@R]7ENNY1Qf
5BEVTXG3&0T]KcdbN_RI^?NOE&OAH6TRYP9>GCOY&..(-4&PH-++^&UGdECW[4+I
?Qd2VC+HLH(LA#J@2;\6<@NNb/3#4gRPK@)T69W\bHV;G(4[JcHEbJE3bbWX9U=,
=?NP3N\;Gc;QdXd=VY<VDcKT_ADQ.5@+OB<32\bY>dS0U:3dJ?TH(UTB>33AK,c)
ME#:B0JaKg,&e/67]5MK.J9V]P6O5HMKc&VRS-7Q:<U2U]>NT^Y&<G140aZ@P:cF
A0BA3FXY30dDF6THKf8Mfd(VVG8fP,58Z4LS&g:H?cB[N]R/4QZYNP//7=BTJ+E^
>-^G5JEX=CB5TSLZ?@Pfeb^TSB+V>\#fN688Z_2OF[eW(.^==X##deHP:/;gEO3?
)W#H)-e;,74<-&R6@O[ZK6PPI[NBa;/FAY004#Cg]7G6a_/^W91AJgVg\?XH(dL9
[/ZV/849MLA>4^c41)#g.U#IZ15F/[?+I7W,?H#MKPNdDN6^,dEG9@,-.CbaWL,Z
:.+-2[++g,bQ)3;N_:TcL0[e:TA[e5JS6/YHCUX+X/T_Q+Ef?b=&K,@DI[HPMaD/
O3Z.a6;RPW,23d@N(085:BAf&c6?gJ1_GZAb2MDDZJfgQL7:G[.Q33?dCOFBQV-K
2]<@_cTC_2WM3#^^e6F3<fJKMD,824QPRC5S\U-,K)W0[18/,(TbUUK2S-BNCaT9
gLD_7\<JQTOXT/&#\Xaa^291[/P_&4WdMecJf@RB4I7UY-]F4T;HAQ:,FdKdM)R0
W>0e<;ZP@JfS6D[/W1>H9c,g^1:6TI-[3=f-GUSKMa3(6<66DGPYJMC;3X]Q+8B1
>,b3MgP^0U5Lf?])1@74bL@_1VM43[ACB->X4_Y[P#.UbA.@YW-Q.Z)DUUVPe=CL
5P55?H.)C,-]c&#E(>dZ597O,J\Z#c,30ICNO;>_cDB>aH:U#>9ab?P2BGc8I\3:
0U+LaC4J5+/_\L7,:DQ2C\^OFNbP,)0@)E@Z+Y3]Q:P#U>:-YL3TRJ3HIg8#T4fT
?(5TP2Qe8=f\M;dDZd^H1BZ2_DZQXFAQ.>>S?#H1PZOAA\F0TA03;0;Q6_3+;YT\
a_N+=)Kc0D5,WWK5_HbHKPg6aU9#GRY:)8N-3=8]&4.>._4PE5\^_]9\Sb=S>D<Q
(=H1F@E40OMAQTW-[HZ=SMN1\&I><(:L>MQ5#.S;B=&[>#6gZEQLGPEc1JO/gC-#
7S5Q0D7QZaC;U8d0P[=W:UWM7M.G<3Z[)QWf);XT0gTDM2TW27J52Z>aL<63YM?_
PZHXOea]M#UScZC@[G)77LB1P=#Kb7d0Y;O\LP?KUSQ]7;@T.4XJLYB0JUDB2NA3
?6Mg7eD[&aVQ,fOc]gPUU<9Y2/,:bP2Z]B0EGJN)3d1f(<.&@A]4@1fTeXOZ28+M
WfOCMWBO2#A-&BD(.Y#ZFLVFQeM^f&)Ue<e,1;-9M8U#g9(\5\Ba40@S920U1]XL
FQM/?gO<K4g])H27-T/FCR(8)9Z#H5CPA3Y[&^_G(S]6MG9MeBGL_8IK+IKQYW2.
UVc:[<VDLD3M^cC24.G[f<PXKWYG8(]c\3b(>1]#-3U#5;BN[((L@b2MZ\)5gY)+
DCN1Q5@U^[3/Ga=RR2=b[J;X4(VRfE)=RLM>,LLI+56\HW8H)AZ[2gEA@-:4A\,I
>QYG&8Sfec:6X.N9K9UDD2Q1)DMY3aEf9:3c,^:>E?E=0TUB+@37B+eZca,DCL7[
Z/AKdEZdIG?f1a<KbdP.NW;R&NF5_PL3X21J.d6[GGNHgcb^&C&[Pa73-1]PbH_R
UZ8X##7,^>(?R6bd</cLYKcW3eAg5F/Y9ARf_4-GBMf\eS61;1Ic7/bO8\c\e=V)
X2=J32Q.#EYd4M-927T>1:8O7+U3J/[O,GJV?F,SMXe@/PcDE?f3L;XD4G^O9b:2
7^EfJRH<D7=((),>\4+1Ua4[]5;]<eRIcTCbKZcXIX+G/>;L7cGJd9DKQO6f>G\,
4d.^Z13FM8KMd1A&\6?gXB_(VTPf<#0XAab9aCFBeK#7KBTGSCc_\)_7(KaHdN9,
W74-LGB16XdO4[-(V5.]&8:71FMZS1Q.5==NZ8b>?AM_NeFEH3Kb=g3#aRX5=G0U
Y\+<5RB=X_Fg36(Q8^/3._[Qd;95e#2g-/WFD\cUP-TcX4XgT)_PZ[/(4OY>@U77
9FTPQX-6?.7/YO>@KN79<c.Y@eGTUYc]@VKa\M))>P/,R4.b&3N4)[g2<9cNVQQH
;O6-5g,9XZUY-;O@1V>7<=bYB>#G3MIE?&&VdIKfFG&Y6?.Q(BJ3VL6=?GAQ//ff
M)W4Sa&0AeQd<Fb]4+(8.4.?4V?_RQMVHD;B2e_J;:T-U6GVe.VC\dP[[E(ScQ#H
SQBD0a2==8K)Y:005e++LL_+F-R?H\Hb]8)X59;&WEfbg3YN_T5H0>-QCc3H\@V\
[[(3M_?@?eM81M>Eb.[K25+HWg)9Sf[:f>/M&eA_)fU:J_/:UEBe+:gED=V<ZJDH
\HCL4&B:P)Y^,@@\2_JD0..EN3A]+a<Q_T&I)[0@A?HNT5\P(<BZcD@UEaVJg+gC
dJaW6T3:E7FeS4WV;QH,M14+0N7F7-OcgG,Q964)WX3[HT>Le:@-HW&a/9UP_GNH
A@[1IOE,22=dDdg,WN<&ON+V=0\a\SDR\R?5C:B.A5:&4>:gPC6E@#)HOO#FWa&Z
)1JI45228C,Ea0CT-B>CCae)EA(>GF;1?,<,VQ</S3aE+749XOWAG:7QM1VGMV^Y
=J&cCb[(-_Vg=E+C<[V]abcg1J8b,/=7#Y2DM&\&&V@C^:d@@1ZU_E;#C\KLHBeA
WR8\HbYVU0#R[5HG;2bE6Y7P\YAS<gUH:?2<+PT6+;WdM85a0+XH2GY6\MDMaIET
3]J&aB8aDI>g1g0(#K96g<gS]+5R=R3#>E=,#?Y5WD0K(dO4AZd&aHaM,&ZA.&00
Q#P?eS-IaE,8bS6-eD9UGK]BRL=2?TPgc(F;Z\,[@gbGf)IUXZa>e(:FKOD/P=,.
V.B^T=8:VOCGQ&e2J17URd6_M^AaOOXA9Q[-OUX.a;HR6@5bTNdLT&;CV;?J],A_
=PDbHdW&aK2PI\(M4L<5O[>@2SCB_F2>eA?H9VNbMK,JTSEK7;2DS6OF;\NcFVT0
#Y=eC>7P(Ua<X@GT<B4HVgQW/6C]A:5-Da^S\\@aR9V\H_^E71Ge<WRN]#GWZB4c
LJE6XZY.eT1P+f+?F-08LSA./\_L6C_=S6#2a?FKT[.@^582BAE8FKP2,fL.PY?Z
B-c7(C,cP3ZP7-@+cL+H,2BP9SdD)L&U=8e:Z1D=]cNX7L]FAbWY>^Hc6A@<N)&\
Caa,:DB@>8;(R.,cPJQ4N:4OfIbd>[Z?2/3CFHIN2H2(Ma4P+JDL1@c(21Q)OU@J
.)S0(afT)EYGT@f08QPRbMFD>3=.FdM<FBV.We[EWRB\B\cMT9QM(5@Y>N(U;fTf
FF@U2R019/fP/@;BLPDab#;JaMOYV2I0:a,;DJ>[K\H[MJdO0+)F(&V/BO1A8PF@
&HJSF[dI7-JY2FGS^U@RRQO6a]LD,A<QBKP=6]XP,+g,MY.H2XE^WV6S6ZQ&\e;V
aPeDSV]O#L>F9E+da=L,@<N=1@@b@/YC071aA44O3bC=GCFP>TY1[L(,&B[Db(]<
7-;09S;#W=ff,?QJ2>8VV(cR82KJ?(HQe@QW^SXF?>9M8Z;M;RHQ.\@_AM+JV4f[
PHPWDdV43JZ5RY=(S1=FD04Z)-QWWKZZ?_8(4c>,_U@_;=L</]^KA#]JSEC9E4BH
)S<U]15KHdD\ON?C7><IHCdE_^=a;X=+1QP_U_^e,+6GTDHLH(0[M<8AZEA?cS\H
WG:[4M(5)IH@f>@H4EfZba>e@J0BO-FVT]6KH0=#dO?P4O3#@-XY\U+NZ,:Q-@B>
(?^8@dG,UJL#PE[gZH+<_PJBc#+5Ia8^aQ_483#XWL4Je_HATCWXH5BWb;\GJA<\
2W@HUZ@bF[50=T?R\/+-7F\6cNH3D.77OO&]75dE@//YE)a&E&[@&:Z]]X[4]HX+
e,c-cJ#0+c9Y6WHJW.I<T67I=ED,29R>V,H:c0g,N&Z5II:)=J<BJ-9\)R=g5L_C
M+#]I<C0-/5EFJA7FaN]0IJ#K?G3)1D_^fdH#FROb.963d)6MICJ<BYL;.7NLD]M
YL<.&Wb(b]67/#[a(-.D=b0N/f4BgJ/fA5<#91^VZ2T70Y\.\D6M)-,.B#5:_4H8
P:8:H^=Z=C#;H5D28/Q;9#aOg0#U\T2U9f4V>9[^I\V)\>f&()E6+:\R@c<=3d:e
<?KSdc;OA@5C2ONO6K&be&W>gSd20DUaIeIE_NIGe>[XELO2V?89^\6]eS3FbEZ4
ZbFN3PT9/F5>F:9/1[U.[CQQ<PRU7)@]U@Z#?3/RCcdI\E;FP>TW&[4<&a,,/5/^
XS-S9LZ1M:g0U4d:feK)cc4)43aT@e??AW/1f8;2@>?2+W[>67>JG0Z3DF1-fL3W
g#OFIY<_9R1bfdXYb98J6H)4V#^@0B71L:,fGQD_.S=V^H;:8\H2)99IKJ.gCJ7]
E/g8aMgU+CcGaF1_22[L#WVB9)DFb#7(_#:a@W?RGa=PYTNa-+VX3;,O^RIG8O:N
]cWF=;.ZD>Y;[/RJ@39+6(7NdV=L[M4F?=F6-P)K;fX#GB[gW[9XD8f>/J@BgWRJ
VOX)cG&+50L<<-b6:H;_[3AbTcT<:549UXG++_<[PPc6L7TdS/P#6>;QW0)Ya;fK
RF;[=@@YSK?B-CXY[ZQg9D0HRE)/1R.)WJHP;J#HG0]U@V.U9-Z5XDd,(BD&E8@A
:H9-NeU2VgS7d4N3[ISE;DbP8B,f3C=@4[<C2NZY]1dS9B8,GFcQ4D>E4JMWH;T.
6BQFG^6.2>/\>6TWa-7_f^V#I/8GbZa,M&fa]^.DJ/-O[)O]&-0<---Ag2._3&C6
_:P>34,1^(B[4W8R;Ld];.7O@/6IE7:eC)H&7b\g#g^dNMd2g)LNPK52<JLRb<-)
f5[5?[+K>:4+)b61\51Kd-)MVV3.6b(D7=64]aF>d[?](7V@dCVO3DcOa&aZU-&g
-_]O>:0BK6B)A8FcD7O(Q,.KU_-)_Jg#NH?8T2;[f]XeWVcQHB)S<#W0dY-W2Y6E
V4eRWAg4+NH6MM(2[[<VgTS(XH;J>)J2W=MF?B#OS0AN+^,ME4O1c0>OF?GW0bQ)
Ea:L.P[;;D<@X]d8IP^TVJ.,?23>^KaIECU@>3-DYP[Xg)>)_<[WCL<a]Z;3eLc8
?+VB6V8J)JHJ-<=5KI&5-FVR6fKA-VI^3),703ZPW^.f#(O^)RDMEcTQf8ZYF8V+
4F9?&/>,d<dXT@72RIf(Xg:19Ab0H.F&((D&KC5A>1((.XSV@BcQe:S@JL=;+<#f
:>21EA+M2#NZ<;5TFF:2(A2)cQ:(C1<42G/EB>UG++57d?DQ:H\.LI6+TdJ0g;^A
YIF3a(OU8--R\P4IM?ULUS?cWYg=2-?X+B8&V^RfC-PV=f6g,/.C0FHBM#JTBU+K
IEXb5]b>SW+V)/._X8(RCcD0O47LfC[Q4f/3B2eHHNT:IbA[FJRSg4K8GQBK&ZSc
e/>RLO1&JR:6P@Eg1F4+gV<eHH2FSY?E>b1/P^<Y&4</SF365#2O/f^>?;eP92;.
^c2HE&@AIUdb\0N]UN=_^[K&G9Tb=C;&P4:_TMW+=WZ6Ng0P>[>&8WOC-5KN)5MZ
7debC[8>#1+>2S6658?8P9BABaH]=?Zd26e_gKBSVUXOTRVYIb9\0]_R#)MC=]gY
.I?dH#dN4#?DQI\6G3a7CfJ+J5:.2][S7@7U7?OdOC7=-)X_^HIOI;&Q<H6a@-/V
+3:N5e=K)XH-R+A95(e<=,)fK=]2aVM=]7+5B^aUUeeQ=PeU_#2;_=0b.OAGeVYT
_e;^CQ3#0eVAGE8Y-TT3NPOY;YSO6:gJ=LaaeT_#Z95U8gPb/#8bHT;@&GfKP#59
7^-)f]CF(fZ@5(CBG7RX;Z4FN@;)RH>f.DbP&4;.V\O_H;bgWEefO?UZ_969PJ],
a6?MPM)../X;_@J>-23C?FL2Z<P;P:^[+?KJ6d4]7&1[LL;H?.cK4cbbY(.7SPgc
ZEWE=fKC5g#/GTZB?;Agd?FIKd108@RR].6Ze^-Sg+.F6@dB\&/N;-Cd8S^KK+<8
LQ.]4RX+YKLK?XLe;4[5<Dd_Y8LA)@B4DU+U]P;3J]W&&_2PD-8Q#+4\54f/G]\c
;a9&X@=5fB@b19F2^.OK7]13CO(5#-fHI7PaW_C@O7/@.S6Y?Qg<NF3\QVYC\fP6
56/F>-V07GN<7=_/3d,7Y2E0HcD?>5^31P1d4Y4D9Ad_0Z0Z9,e+B(XIUKNR4YLg
]ec]:@g)DE.UaAgX2F3T41U;e(OgPaISN7ECcI5GOf(ZMN0;T^/9b8@,6/44Qda8
XCO,_-@AIG&4#D]F>@:Eb0];BbB;WP0DWUO&;W=:cA4^fW#/V16KSH=5W)SY\0TI
KK,gG/G3Dd_>8#]:7@IF(O?4@B9S[f:,QP^de_E&RQ/D=KIZaFV47,\@6AJ.]P9f
@/6M(\90N]7=;fb0b/)BNAY&^;:U42,=R#[A?0D)f;G+fa4-X]?=Gb571:VDHH/(
3)#3Z-05&62I9=O#0^.Q4?MY^;D1;MOBPT7cf\K-@YL:0]>:#gH(@0E\I[e]S&CF
Y0]<BJAIK>4YN)B(YcR5HA=Q(e<HB+<>\-FBW;KbS^UWWg.:cN;E[SKX(c\AGMKH
3B),^\D,C#RO?1T=Y1D=N^W,GLFI4V8GYU6W1C2Y60I1I^O2[Y&1[&>]>-94NP27
9J,=g\YRBFO<I94bG+UD?=>.U)-(B7,e,?]/NB@;\PA<-KM;E9.#7+IWC)FU+\/O
X;L_RR-gZ88;,Gg-+\]I>4.7Q_]0Ze8-M#LX&=M1JY4R9HeP-IYR.-:]O07-7dWd
>OH[TXQ,=<&Y7f+>-(&d&H5\80a39E32X+,0G\S+e<#Oa:+M6DKgDYLQ<Jg5EL=T
_)Y\+CSG0I^7XCB?SC>dU]Ob_-:86@gC2V8MI4)CaZVc+]MVUP=3U(DG0=@B=^[f
IO=N&HcQP4G(QF4++NOf)#LWW1a4-:])&G&+6#?,M:82?0VM<-)[./V@EG2^P7/3
J74b5)Ve8@#S6)X23-cHCCgZ\OY)BaM(d^]3.6X/1O^_B6[2QDMaKPUO:C0LPa4[
8(QcPCN:_&)Y+I\g@cZb;O0+Y+HF^^GE?e6<^I^\JfMGN^73,966AdbV4MD(<IN4
,^4,g1B_0#>:?Q74.3ESC[YCfR]]WT2EOQ7+MVM4>\dMcaA72GT8;3?&O1fa:@2(
EYU0WeD,Q9:ZQQ5_L;;&aN[,A?]ASg_<8H#&bSMd2KgWIA)dDV0NFgY1.:^J&.-1
=gad5&6Q^5]f^JaI+BW[VeeU?7cLP;d8)Jc+A_(0LOUKRX#-NYZ+GH3]Y/1]GY.(
1;)/X9bQ..M]?+B[]CG,>.10X<Xf#96,()cdW:W;^O@Xc<f76(S4b_ZV)aW45#IB
7Z+6E&E_G2\R/:9)J]FI0?T/[73=6C^Wdg1Kb(O@HJ0>aO8c/F_6;LUfZGaCM#8]
YF/^Y,UB+#EA4G-_4DIa10cFJ>VLJXK_C2&5ceZTN]-(;S]KOPLXAI5,CGHF6@Pb
:WQ)MTc<c7M]87bIdb5_a-^D5^HH/X1ZV6@JB^^N#[9P#0=)\bNN0bV9XX:bX.Yc
>NI\CV)2B-=fIOR5L91a>g-SL.INb?ST0bS+.3f&e@-)=;f#B.>R].WMTTFUQE#g
Ic5B0[g1+Le.305KM\_W^T6c:cg4bgIJ@XY_R8(:U65C,?DH+Q<PH4,)U:8)_RJ(
C5J\TgPHT47?X(6G3-:^b6)MbFc-,#5P3R_U?8B,f2Kc:;]3N?eIV&^JBMZFSR:.
OIcD9R+#daM.E-Q?JdW4a/JVZT]R5,:f3?;B.e=;U?-B,1&J1A^J++OQ6W@g)Z0.
MZDAdKL)K;L>]8cB?N(;>^V(/_CI_-^Oa,:e08Ng6I32:&Ec_=L._8L\2>Pa\\G(
)@QYK]gg:-@JFe&LZE.T,;U9BKISFN<:M0C_W^BR]JX3d/B3a(cO<EXb>7-Z/;:)
=M9WDOZ\YW>fe@b#KYdVRT@PE)IMNSEPG9(HP^f<X?<S3dOKN;CL5/^cbB<KaHgK
f(MefMBILfaY(Z<\EFUA@2G?PALHC9.R_=8:cXO_W(KRWP5a3[X46^G;XZ05X+XN
^^E,ZE0GDeTdd)8JO0+g[#d3QV7.]-</#cZXYRCRY=3R68[+K;Q.3cZ]g_@@@F>d
dP;^4\:-JJJ7AVBV7I#&B70G?[3B6/HZOa?E4OJ44F(&g6\:W-^IV@TKLJLN]GN4
3#\7_/=G.MB+6QKPNLY[L0U?e<efE8[X;US<OO@6V)9N.^X1aE-7^58-,3UH\+d#
N+,]VQ6XSQAD7bX>b/\gL7(LZ.,^[LL_8&g::.2[#M8H,c4cI5GB\]^EBH,He[XH
-_1RR>gN<W\dg8W448(d>>/M^/7(?,cP#g^Zf]T+>\WM>_e:ecY1N?&>M<aMY7<Z
H?NMaBegd5X:@ZAV;2bQ-9S?IXYB-@;f0?fHQc+(VL[>.KbHFD7e,=I[>:6^V28.
]<GZe=b/-BDg6Vab_XSaNa[TaK.<0EBDd;2_7#P_73]N/ATQ.VO;P=#3ZMN&YTVR
1L/Dd?>^[L=BU&G?V\\2E013MW?E,B@&R#/R9+<RbT\=#TfB:4#-.0/?g4\9]Qg@
Te]D2F7(G-P<-cCPA:aIZV6Ua\dY&:1Z#-gb#/KA.GH+6OS/WC:NP(4JPe,fBGP6
FCG^BFF;Z.=V8HF7E.9P,Kg++ccT<@BgLgUdON1;ONe4T:]69a0VDeSK;CO#FS.:
-FOSL5YVJ?N0Q\Z<QMSgREK745=7V3AC_D+Z@LERbe;#6ODgKWKM,IB;2Z)5PV-;
GUSUHPWBM4\ObQ3NM228I>:,#O]H0P_A0Dg0>-cIbKV>>[a+B[7(ZRA6P;&XT8/9
C_([>8.(+DHE[0ZYO,8<0XJUI/9[#_X.2Z5TTK>OFW[?EJ=V^Cf9&EG-S0<BVD78
#6c<fgY33?76^F,bP1S?L4\OO:),Sce>UJdVZV8]cY4UfY_1NSMg)#Da:HGaZVQ<
(CL77DTA@#NcPGYaHg+D\-E&M_XVH#_H<X>)[0_BM^G]JGbGFW>W_)AdG[D^2^7<
<9:)_H.2U?g>8[T@G\fW3I4,AX]1L:LI;BD)T>)K;=_#7]fgAO4\#Z3P);YNFcg:
e43CEdX.6Tf45S-(J8I.8O1J3Sd_[gD-[4X6:93<WBCcF1Zf?OQ<I_Z>&FbVBM-0
;]JYSSG,-<=RaBMe+H;Aa1I9=G?JLN.6g+a9GTeCM)e0VJ;/I@WVB&6X-83XY.9f
_O,D2Jb=O,OEWQ(01EU_C99,<FZDRU9d.^R8NE3gTE@&3+WJ+E,>c#L32?2UZ[aS
_^f5&<86+Cb#1f<KT@b1:FUXPG8F)+8M/:_CCKQBUTMUWTM5Z&M]+CC;R;e(95P[
YN0U+G=/KKR8<_&V3@\32^\(.&19T5\DMYHUaU]RW]:<f\TN(39558P#W9@9+FD2
B-REZg8-eKe@>Qg\)9W49T=T._5[?VR5G3Z\UbZW<X/+LC6\DD@+a8?cVM#CDS/1
+0Z.)7a?P3<3GQ-J;cBF4Uc)>Q\-1P_1K/&.T??^a=A6=6bN_S1B\HKOAG]CL6,d
?M;3ICN_GIXf<g-(?9.(VcN0TO\RI?BW9+BU1A4EB9K1QR0;]WE9HaT_[V37:eF,
T^N@D:_PZ:J7ZEaL>/,]b5A21CE3.@a54f<9\c4g;f7^c=;cZ#HIELA_2VEU_)7;
+g8Rc:H>>_]Pe21M:FW5N+JK0cBa@@/XdW8NDCaLAgKP6<c+<0HDO),+EK^MU^>N
WeQVR:=3N<a60g<>;[?N66/9CXf[>@/e?@)\7XRVVJB5H0fWdOfb<2DG.+8DW@aT
,0<d+EO?1]F,]WAKS6=P0FM&3ROI&TMCNb/,U(J4Q,adH])Qc-SJ7T4\MM^f[f^a
eDUQ3JX)<5A?93I3:MR1C95\ZC+4d_+)bCad2S9F#BHFffB,O?If9R:V=gHFH[a:
dSBO4P9OT#+\RS)D/Z;>1b@b0ZSD>I50EI/e0_.a@5E][\9,TS.9>Hf)9g&3/LJ&
)3R;@/V&B&S]3YLENBa2]S2^E;24LdBWdM_gC^1gU0;5-=[Od7Lb\Fe2a\f07;^P
S4I<0]Yb5B^?)L#^DART,N-C?FfQG#Ha)0KbTQXY.=NfgI:a+b[8V2fLNFKXEU]c
:OC3>)Z4Q]LMb7T<\P](2:LgIZPT[,b?+MB_]+9OS=b\QBf)C4IHdP@(E[Re0eFG
Y5_=b&J)M)b]e5.3N-8)=#JYS3]eQ88QYWO1cNfeF[R;AeML6&>A,:=0LHVg&_[V
?P2G@<Y?c[Z7\CK5]T0+a0UW/)NHaGg1e)>?_E;ab0.O>:b:?Wd-&7+-57df+QXO
>E@K,/^:5.W#<R)4d#(SA:B@&2E.SMAMAEZ-4bM(YB6+=#4BL6QX50)T:2FQS)&2
F?@V1JMeAA867^S3Hc^[Z+A39-IScd?_0H[a?<1OM_:;bDTZK8N8;L)be9cJ.42/
HK3T&H&N>OFCONb-.g(,cQ54TVWTIOXCAV_.VVFCW4gDR^WA4(\b^-R6#&ZJG.b8
1&f2_(+[+KH7N&R@R5K_Y<.ZO5RD7,\;CVe4\a+@UN7[9T=Q03.QER61f?WOZ34)
GaNaLZ(35-PNfG\0].g;P3-;U</,#X-dKK:UHCB<1Af.HHC7JIa+PWE8P19Bg5##
UdQ;9_HMFffK@:MP7>A8ZC;9QFB:,gEF5.@U[<RRJ:cVDb/EX;1cbWf_N.=c5f2Z
L;T&T8Kd/cI[I?PC7_+3^#8,+USK>_2e&d;g\&L?T8EYE=N^K?=\C[H4[-ca?F3G
--5>R<W]bX?F(<NIGZ,/[=922\S3>V6PZ:T99??:->,62]?):#G?_U,>0c9FCQWI
VYfg=9Yd:^0[^,YbfQ)43,[KMK3>IGX@E2E]g/G4Q3AMTXa1;\;Z_b7B5a]bJf-F
5<>&^F^0LI4A+<UF^)-RZVga3IQ=>F>\\RQ\?\.]58C68HX&(WY@63/:B1Fb:=Q\
K::A\XK/W=^e8W>)1@I?6;ZZ<GRIP]=Pd8KTI0&@dPHVE@BLe/b_GV.XO2]d4MBF
GTgaR6\f;c2#U3a2g-]d-@\8UaA@@=W+7:C+J?GYX[X(c;GPe=X&>/\&@cgN05EB
8:,)=JIWOc8ZF_8bf<#@=9M>/\W2</+?1GGGCO4I.C_OX?QXfI1R)WQ+A5G(IgEO
,4[cf?7?)&URZZbZ.KG+0PT3Ac=ABIbWO37fWTUXf_91B6^]@g6(DR6-e8/EA<59
LDg?5NJ8=>&V44O&DZBOV&#_8X#V>-Z.WQH[Y)0#[?0YHeb0/WM7CI0eYY4<\O^M
+R5J[<\8FN??;X#cJcHVWQHd]8:O(D+F)<E(c-+#?]5LD8\;e;5eYYKb@A6GXN4=
\79[[Wd57@;(LJ985KCQ^VfTG#ATBEL_PgLYJ^O=6Z4X1aZJ6.3B/E\1SXa=:L\g
9I2GNHP#M)D.:8W.YN2TV3785&AgS?XGLM[)9LT?U7QJOXf^a=X6\YNX]\7^,DPO
QL]4LF5e@;R#,KJcAS[M4fB:\DK_\-W+0LZ522TJHM-(bfDN].He+=AR4P,?/FMO
&BWa(U:b:@1L]Y)-dd^99:cc,GcP#XgOV&?&:K:RD)1JX.>Ya7eI^+UHRO.TIdgE
4@QK2]P\@[&2UdYcHf+]e,[LfSI#EV](6-S>7;TZ:bQTDK0&b+Qg4NCH>g)OSe5A
4PMTe],D.-?R0fIA1O9R.;Y+8[2,Rc\53BFZDgg>.],SUYLc:/&/^H8OOUAA;We#
Q=_<OaFR]S+_.X[HG9QgED;.W<1Mc^9&fV5/^JBO-@cGYK83;:+c.H5>9I+E.cPJ
[.f:/\4X1MV1F?R.FU=J5Q#c;]V56:7#AXPO]\S\fL]0?7GWEYD8bVHKH/8a55=;
PH)[=A/-WX;5+5U\,JbH2Q=D_(_-dU9>+-Q93c2M0?PQ5B.:R>(A2b4e&JL\W0-^
>EPXeC6#QA@S<4J16A?cb)[YZ0;Ncg1J8H.Z2M7>\M3-MND?:9/J_MH3aaK]N/bS
F\09TZ-..d0GN0eC1ORV)KOBObLN;I#G=#0BC(R\4Q]YgU?ZI+AY7^VWa>UAc?#Q
@4XJG5-+G/gJF37g&Q4B\9B8gY#L(6);^OfcQd&^J3SO08MB/_#4F(]2S)P,:8Q<
aR\gK5^H&SD=D):<:>UbA;&33BTCb-L=:1Q,.Qec3R?/O9<0KXM9RFTC[CG6W)&5
WF<HY@(82,H+:=6IY)9a3YX52(Qb_/7/7(fR[B8;Jf8UQHRAY@NHb1@Z\S5=+]0Y
d6VV@YI.BD>FG5(1_&dXD4QN08L)eH><YT]?BISI(QH\2-DP_MRYHI;=:EBQ?S#E
M@^[_V;\+HP/>GHP1;CVT;0)>J51D</f:9D;Da(0)S-\XL#VaS6AcAP#13JCgcFS
5=3A+IQ4:4NMH69)a^=f,YT>XZH+3OP4?]KPWPf[6EH)YQ@PBM7(D7<V=UT,RZS]
+5(Ra#S:ZG7eZeFPZ&5<_XJZ^e(Q.E@S(^19EFZa]XTLEaCF<B8Me80E)1aA:BUU
(c,0<XG]CD^?[=+Ke#gSe1I2.;,0DM-RQ[[cJdZ<f&d=6,c)VbaD<YX)#F)N_JO)
PPgXZe4:1[fd7M(.#A^>)f21_4?DI-/MMY6C0@bZ//=f=HeZ4<\J6\T?\<f\X&GX
+3>\I22S?P^Ag2XeF]D&P#IZF/,Zd27-3:U,Cf,=DS,OL[3L,=Ja.7.J0-58+>e1
44=HYFD\L3KH(;c#QFe9F?Se=.^6J.>C?:/KU.5EWf.32fC,9RF4>XZZfUC9C6<L
N<?<#5-X70X@6_acJ_1D8E&AF>WQ<^VJH3,S7U4gQ)EEHQb>fHe.R03<F[bFU8RG
1Y#=++b)F@a#,FK(g2>aMI#29TO\Z\d#4-1&<,G8g./9C3LAQY(9gbKP&P;7dF5G
fI[F(_HDaf;Z(-<D[:R7WT6HWFI,[J.#QI4^,aUa9[CPf1R[&eDQ;/]UL)ZYLf>_
F@c0gf=]&[<CDJ>1I+4/VNX@>K2J1#P.?Y-9IOVC[FR/,Yd1?=XL(#&eHY(X@a]N
Sc<<@:T#]V[^QGWEHBZAZKG>V2?;)_4N7d+3Yd^=)BCKCbN\U6I:4[MVf=)PFXJ)
[:)CNM]K6/I^SVS?HV\/#U(Tf?b,>:B,<0W^/248gE-8aSHF@NcK](b[1NfC^=aE
9Q21T/HfJ;XeW7d(M)H+J5#19Y)+&(D#-4fAW+)dGI3)>H>eJ&_NDS3<TPH6K9J6
FeJN9I\2@<)3NSFdEMa01/B>/_ff(DDJF503D=41&VXQ,2)7G95E,XVaM<cKQ,Wg
7^[Cd+RHN86]=Jb4f=Bf+P]I6TaF+BEB=<CffRRQVG=F.SI_E+9K(aGG@3EM\ZZK
/GY6b@g?5M@+-OANJJ\L?6Z\d&>\/QD@-(V?FC9b?3_ca3g:=;H\YbGED=[#&P2Q
>HNeLbJFQZeC3(26_5AFQZC8)Qda;H[gW6]Xce^HI_]D6JDZBIQ60b;U-P:fD4K&
JH8F.1<G^9<fAD7NFfJ?Z:b[5VL#S3YY=W&aO0#.[_KV8c#S>O-FPBL>54e=Cfc(
IDW:C\Z9NW\)OF,@IbQ_#\5.&b_\]0,JG\2bR_LXX\2I/Eb)[Ia3MM/R2#R2-XH(
(3:dY#]99(CV[&(Y9YbTdC@/N;cb].^LU=POfRFG?=KU&-\HAN@EIS/U_,<Af9K+
C3c43R:F@LQ<]#APEKDfUK7NAd13Eg4SI#gLC4&=Ge(@/+I<IS=>g:eE:bJ^&.=#
_(9dG.B;cWA&#(GMV?K\B>5L/&[d8>99a)THZ2;+X,bOD&#;IRD[M:X;D@T[62OI
TYNR)IXWe@Z#/B>,Z5;=B4UEbDEZKgC#:QK@e&O:fe(#c@UT+7fM0\?A>/d3#Z/8
,H(a\>V262C,MG>>7@eIdAS5-F]6MKce9C/Fg36[=KL#-]fD<Q04MY\:d.A<_JcA
aC3-A=eCFUDFD.>A\<>G@B4eAcfOg5I/-f-WICd,0/eA?=9g5CW6-(.e71,LA#Ld
P/d/aeG1?,F#7Uf-=>Z.,FJOBgKZ_ZM>4=gN)818L:Zedf0N2L+EA6e-KC6V:52[
3.E._J\e[TTf.IS6A]FESFP\R.8@-8;&VVLb+[3?Fc5PU/G-65D@\T+1A0[/FX16
@&TQ?2&A=(d91@[H&H7=?HH0&YEK3V49519\:d_M@N\CRa@&;KE4>@D&H3DFXAMZ
#M&VCNM^AV@e^Ja1bE7X&=#[:(QL0W:RBH8#);\>f8X2@1>PaQ=Z9O)&YFe-LVWD
R#6Kb,T,R6=NW)1;@(YO<.P9dJWBXf9(+-+fTFJYF9?-66&\g.J.UCYX[,MfFWe^
W#IOI:E2+EX8EDI>VF#Gd]WB53]1^<W;/V+SXUEUF(Kd5#4T&-V((c,VZFLQ#_eF
IJ/91M?->J&GaP69Lb4^+KR:PeXQe&:7O>JXVRd,.E&FTIU:6-W>-](MTZ+eJ:Zf
4N9RaVE3cb^;B,<e^DE1L5bM>G<R#R8JU]/_-29.B/(dGF0JKJ:5#<_BQdTcWfV#
B<:c5Z3Nfg&.CYWR;QW.>D37[6)X0)?Zd+GgL-fHJHeKRC6]#TfI?<J>K6T:O>;3
N?<TGUC4DT[),.QF?SPfY6P]\9WS-?;]?(8X[afbFGS^E.fAXX,.<;(5>PVW^8_B
^7UHg/8VWg90JHH(W1WOM,G(U4:.bOLCWe)/GT=B(@W5[2LB&7X4Z(8FMB]S3KD2
\f3aXRPSS7I)N.=.8fC#9=cHYMSN12H9^RAO5D&?3BK:W8>;?6f=XeZ81^A\96g/
AFd9N_]YW4WK60K-F9fbF)aWIfOBE/Ea81d:@ZXN4DOVGZ^O0^SNBb&:R5\8+fN[
A4:Q-U]QEUR-IC9^8GTbP1EeY,\EM[]4AVR7cBN2CC/A3#SRaCb0U3\XMMZH^QU_
&WB3W)QL)]c)TONS]6>7K6C#bG?PR0Ie34K(KUW^36#MRfVXK;\8B#T_>#-;TX0g
d0@f(Y.+:Z16T&ge<54QWS7G;cM@@BMbG6DUMM?-bc<b-3YX[8TWRG[&J_5aN5N+
AO,H(Y+I(J_E21),[U>ZB<HcU_O:/bcV4XDY/OcI>(eGC0\+>0ATf2)4=Ee>Q&PX
gOU<.N.6.D0aS[]NLL-gX6PUd49<=W9TM?Pg=H[3RW9N.:U7LZMfAd:+(CK]_:4.
3:ZJ,<(V@4MU9JJSN>gCe[aK.^5BJU^&X^-2d)VUJB=4b2/G>FAH)NW.c/8S2,]6
ZMb/&Z:f=Vg&<]AQc_-TXAbQM31[bGOfGU/E^f00<)ZE9^VgL9_).GG<A/.<#^>;
Z]R:BW.-L@/86<-aD__MLPNYSW^c@LBTP#NfAE=0P_W.93>Q(1JK,6;8YX:U-9ge
8aL89HO^/+ME]9ICD6L9A.0c+J0]O>)CA8b>;FO;I>TOU^IKPBW]EHLce6LO7.a_
<5#PB0(5<4RHDL1cQ&RDg30bJ,Df_T\WWb1+3f[2VT.Rf6<61IT7THJ&d]]B]cd1
-SJ]2:f[)3,Fa-GbRCQL,3Z4Le/bf:8.K<](bf6^LdQTTP>ZDE9IDZ3@C;dKW2BI
OS+#[WaGOQ)?4QTg6.F:T0:B#QcGA[d;74P]YCE2BNJDR^[MN#E&@d_G^@a7P:.F
e8]eBTMJEWF0P9\88W(8]QA1:S@CVI3be2-B0[[VG#Ng&R68-G^_ad,HMV,[I;3L
Q7B_]GK&E40X;6X5K?ZYGa_XLAa<M\&a;:Yg5DJY6+([PgC&MQa)A_8d5_LO9FDa
4.,FeZ.dHMV/@\HAHEINMUT+@@ZH>;\XVI\aTN/.L,QX1N<T<KL67(]T^+L?(5,0
FKU,HXdGa&_UVXIC[GMT)?3g([[c(M3Z6(g#UHf:A:TX<AD7,KBA4XaM+=>Z(AcY
eD\#S&U^:13&SP03,C)+Eb@0,_K8X]L(R6N)LZ\bT58NH6<LN?3f@/.cdX.NEF9c
_])<fK/,8VZ8J..G074MGV]#5R=beFY3F6<OI]:>77T/JA.IS_:[5P]IA(\G1)e^
;M]c/DUW0dc=\IEDd4cRL;;W85H1Z5H@-e,ebG+Y&dQ6#,.cUSXg>BU_6W=7Q;<W
SH9c62RS:W6-31&<R+@LD6]aYO>4f6O7H(<1fDd]GQg[?L1:L?5H#@]7cXe9+dOC
6+NCS;gO1L+4K_VX2cOX:/[RZ-+BIKLNH#^YU#DPYJK3Q;7[&J_)CbM5RDCJ8JK-
Z3@1R^)NJ=SWRd5EWK;/G;-VSYG=YfLVG1Z=\EgN3J.0ce]+&&7VRCfDNd+LP.1[
20;\NEf4QQ\f1L;:ZCZ]R=VC1N<(8<8YBF-1,)DDWE?^D0P5Vd2;=ZcXgPTM460Z
B>(H__PQfUT4I5BD5F1aYaegVWD(_DIZb-G+QE_B8+2TdV+<[WZ9-+HA_d=BB4;.
3La0/eC>[&e<#DE0:Y;?e69gIeYA@_-ZCA[V@=5M=712?2Cb9^f84J+CHFWaIE)\
dI<6O<B^AWK70N-A@(cHH7a<IP(7KbeaBI>J7:dcM)=/d.WU=H+cZ.YD7I=--VW?
U66F:>Ve,T)NdL5c0_Y^3=FXH-_O^bW8BKUK7QCNcEgKXFR>B=MZOU;VP/G?g0f/
W2Ye/BIcQ]@4<d?c?,E4D\fG\;-8\IIa0.]MNHd&c\:3(09TW^fNG)QF:N@R[N,?
?>+dF,fVD\.7>/@.?&34DVfE[1XcY@<<_XfC06VeYUHKE15A#\/TfADO\aGMd;[B
D?FM.eT5_SD_W4];=f1^e&;T5-64e-96TLR<2=f)?P<K7bcGFLaWNQJA6W/ReH>A
fLK+e,ZM,5U@PTc81XDbccU-NZg+Ue^cD1>ffAEFSF1FI=CVdg?@N(LCHW^cZ^.&
&YR-]//b#L72?9,KgA0Rg0=OE)ZCHHSV09QES)E>1f73386#^LD\4=a<?=]5<FG:
:UXN@[LKSaMATT\=4TNUPRE)A),<9VHGH5OUWeC<3FbG?.4E#DGGeDZc=323?HI2
LFS07;P7<7cE[8Ode6]cGd;1<.6JCSM;3b4(.NELIBL]Q<UBB>C,P>a,Kb<TG=Cg
Z[JeAFf9F(HYaM/?^3gBB\/IeJ5>^I:>58^bD&G6EWP<bNC(.b538ER>cYc#g4?/
W8^=4/6.RP(#ZFZ=AZXK0GTUcag5bIR_?#UYQ@M(5QMIV+]?R[fDbcH;WO5;G0L,
dcVe)39BTTGE5e1B1bcG+\YbJRK19,AGEXK1bK&I^)G^3>PQWP[MBe@,J2J0=I5G
UV3?PC8PWG.6[/IfK73,f.bW--[?c=Q1D0(=HcG4ccN-DU)+:R3S#Ga.@8K.Fb1P
?Z/OPb:YXE/)ZeUNfP(fPH<B]+]_>g:P0V;CP>@5JNEK?>-c36@[DA-+WT]:1@OI
LPZ)KBQDT9_YBI<c&S]PXE7@V=7]_.B[5S@G9VLN8VLg32;XK@ST@T,U->1I,F1Y
A0@[WJ.5-ONHEDe&UcZX.X+?EX7e,24G/;-=cA\WgeGWLeT:G#^DHMBKN]>>d@A7
1LYXN#S[F_EBP&NSHRg3:e8QT0+B3I.IgF/gLcZD97K\N)9.EE)D.<&509V[2#@D
b0&^4A(I>1-I.)PQg(/c&.Tg./,7c)6P#Vd/(^)Ac1GN^W)=+H=\V4Be&K>A+=CO
2D/RS<C.>c,8gQYV@21]YF<.#+KdB#.H_52fNFbf7?e9#TQY@c.Qg@SRY0dYFgU[
B1N_-HFeVRAU8b2?..4ICA=H;K0#+NCBa4d\fH_I9b#33/.DQ36^<F<II5N>?U<b
WZC[6T-BYOK/_,V@LC,0U\d,(KcU,T,IXH,B?-QB80:,M#,JCC;c/g.7S2EF3dU.
IRG])JId8Ea;33CBC[d,KD6=(I0@)]eg)@O2O9NJOQ3(a?@4;YK0:?]dCEe(X8G/
)LILVHHFaVbO5:VX4Y,0HZX<ZP#PI?eUG7g@SeJ90\7&[R.DJW-I,6PUJNQ^G7:,
-,K2a:8K/=M;>E3)23^@+&K@9dQ?[/KSU<#[fXGC6^Ff>SUY-(I)MW6?==>&8K,@
[I=+>_/Nb4#P-3G9(TZTQ;[O?J[6gE+;KR^+S5E#:TXXg:(b-8A=J5ZdSCF_Pe#7
a,^779BLU57=^G@L)7fH,/aYD&;6;G2fU=M+YPYT(7QBYMF]E&LJ,FSc&@]EE,_D
TfB]eA3R@G/SZ(+cf8<T=7XYGKC7b&R2aF6\>BH,Ee/F9X.+G>;=ZE,9bZ=Fb77e
NLf[.1T-7H?M3.?DF1VR?5ORPC?>>Sb@JcSR_,T]KU<dfZH\V6RFdeaL;J:,96&O
0ZYH8Y)^Y6IA4WVE6/F^@EJES,V/CgX(I1I0a+0Ib250ITd98Dd^FKIH3]2N_Q>2
a&bT0R.d;1O_FH5YOd84M?AgKCH#5];ONRKVScI-a\]0?/+c]F)&2J.CfRD_8^eR
Q?&S@.Z:IG,.ZD0BWQ27eU-[1Q0^@+3\M\):I6PX&B7=\PN_+NCY2IPOROdE,XB_
U#b88Z1EFe2M_B:Rb=+]<X3:A8A68E3.+Lg=01A0O6Wd/&.c0(+aU:0X04+1V]73
O9c,KS2#6_JEM5BE;>ROY7&KNL<5]2.O+;=UXG0GZdN@6BKQ/^(]\H^)L\QeV\E4
e[9CN+eG>D=.P+.H@?XVED_KU=U3>:cRUVKdD2YCN;=KZ9<23XZH?dXT-,9CbV^a
:ENH)7/+aITW&Y&/Dg-,1XJQ.[5+TcgCAfI0_7(WgE<]5C#THRHH5#BW-&HB6E\g
?_[]<&H0QYaOJ8A,7:R>?2ACU,g=\=T&P/8/M#,f,BgOKPB1ca9QO#&@1L98\:.c
NCELe,=e>+09^T,^QN<f#&J_BC^M[LN?ggG<ATZ<e(.T8B:eC]7/?YYWA15@6J.S
0EWQH\+&XUR+J]Yf,0-=9+B2_LeC#^)]CQM1QD(#FF-e2#,(S#ECZ-LFWC0Q5^8G
Z.6dMbYYg-6T@GF;+2THF<N]EWTYF0)45>BfPHW&VIf>M9fH.-)=:[G_POR9]3[/
)9:gN65HPM]D/>HI#BE#[8;K6^Z&XA6+B9=+M@=9RU4^XKPF^AQ4M\/(a+3NH8>5
E<\3<@;K^059B,07O\D^6++SgV&@]N_,6a(W2G]KQ-CP[Ugf\92-^.cf_PCC820U
.E@8?&b-W6WE6Vg3GPUQEAbCb=]_>#C?2<I#.<WLVA(EWMBZ9V:-9+0(+L.-cVSX
B]HKP@A#WWD5g\)J4_]0_S<UQ=9KRX+?+\-03/=:a<U>:R7f7Se2/I_ff3Tba_U#
B#RSD<HCP#(3FW(^LO<d(C/eR64/QKYFXL:PLe1Za464eW5-L>T^?.((5JS##X2D
QR^@MK?C7ce_XUV83g\5[H/0NJ]17U:IIT&RNKEPGM-X>RAK_\R5>TL=B&GD,Ca=
FF2-cL+UU:H?f5.Jb1?6\Ce(d[MXXNb2aF+_/76XCD1CeYF)Q+3^ggfJ@0bI8.Z8
1?@]DR+)8[>#HPKLfKV:<>F;7<61f;2,d^8^T)^QPS[#UOZL-\eK1A)P;3OW,4/>
ZUU=7512W4D=acFAE6=Mde#PdZYM,:Xg&dFTA>cU+F@=)<._]efBa4&HQ>/9f&5<
-F_#a;DA3_LA<O=JdL9Ab7Q<IIW3LbN3b=5=G;8HWG_06O_I[-NHWcM1I2b:QJA0
Fe(6\Q]/WVQ9;a=D=Ca^^D(J:3HL[:d-8T,DA0CLUAH:F/#X8T258U&gG0e3?3F7
(_)?#ff+agL8Nb]4XKX6\Td99C6G.[PXdaSFcZC-R-d5S)#UCF0FC[\@4A8RLKS+
e_51+WaI/[;C1\0XS=IVKWdPL,<DN/H-N+]a4J)c(\g.RRba5?(,(J]4(=#NKeP)
dBVUbL#]14:4Dd/?D3V.9If/5W4HQ]MaL-+5K&JcANI\\CYWc:-\He_]\HbKG,\>
/-d=H((D[?6E?.(KO2SGf_+d5gL<)2@Ec7SA1d(,e-:U-.^#BQB@9/]I[G-COYUS
7Ue(9H:WGa[<d/J?.?W@\:WYT35;CI5A+Q,EE>+M0.Z]M(]I<FeCN7/;?CFZeBe:
T(,K]f(HF@D@T)\H28,FcE[6f7BG8/])b+HE2&>g4LO=ENM7>T5f[,DIgK8E3ULE
5d1RDQBN7J]5FgLga3-dc.fcJC[BQ]PDF0F6C<UbGOa60-Q.#X&&N[(]XJK;.I8=
(XD.JO^9eb2NYcWacc5?E_JY,8<Y>?<W_+3)/E#5I/\=X]+4H]0TEfPb5eCI,73d
/:5G?M9##QMT6_DXBU.6V;A@7:92O_\QR^EfNFd^#D80(J?<+NdYU9;-92;(aBU9
42YI8YPAU-9.Q&VO0PG[AVNPYb&:fMG/^+;,?C0\68P6#XXO4(L?6(O.I<fNZ&V1
F+g2_Ha>g)DXE>O,-[ffEVbGg];W1/LUGa9JZ:6,1_=B.VBONNdeR;70U;IM0b;.
NB+<[d5MOM2WSe-bH4I,=KVNOCH?B,BRA8Rf=d\2Y0NJaU;&K1))RT+Q/8,V7:BI
.G=<OM86cHP(d&\Y2U),5I\_MZD+M8BI^3.RHa<3\7DGR81L#DZP3GFK1P)5M?.T
[H>:d_4-0RN_4(VO5T=[H@3H5H^1?Q_)F-AJ@_BAW-\9N1]0dWRO+LUVK1U.94H+
6c.-(>e[P72T@7\W^(;]8aQ+Z71>-d,ce(WHeA?RN#ONR<YDdE#T,__>.VFA)OB?
SZ89b/U/HDNYAPgUF7:N(D0e>g=L:c>,V4S>)c.)AeGf4KWb9MXIH7=f7?AI0TF1
;W5F9fN@^F8ZG\T22#9:/GD3XAU)<5ULT(3/H(SFW/,d)IT>5)]I\?ga5:KE_.^]
R_VVSOQbFaBJ1)1+c-R&XgY4V+=O)[(+2-TM[SZ@SE]#aDMaDB\3b@]T\6@?:+Sa
-EROKWY2cB.BbE/cNUJaTSH4GK)\OBP&N\+TDBR5dGS,?\Y#([8Y-AX-H(8I^g=H
E(;1MIQH\aQE3b@_#D:^^[QM;5gGXg\g#5gEC^@=1]E#:6M#+C_4AQ&(J636c7P7
b\5+&VU2O&N1VKKKJ1W^B^\U8+]EW/JYBR-HLTR#,JIe[OLC+15;HSA&@a]GFPM?
8bNG88?WVDBgC+YE+B@C\\JfZ1>b=C/4]eXM/M1g6dPOgf&]GdZK3#Obd4&^87Db
,)C<[+8ER3=2(H\(0d0@JAXI73AR-5<Nc7L4:RQQVYX@Q3EF0@Q_[91ZG91U1cRO
SdWJO1(d2#;YP(B@D3&V48?&:[eF8VO<<<c(PfHL6Y3I:+FLCF=-9\K/T:9M3WX<
fD#e:]NP0^A;J2Q1-cCO^4FT^9IQOCgN)RUNG_/NYd2ZNWO@>(#C3_S#5)cJ28RA
KB4]0L3^?Cf+&bd#(9Y9FQf2)030L-N?g[#2@UJ0+VPd,3(E5J+/Z>S@P[e4bK>X
MC4]F2^c5)UTYdXV#7ED-S:061FRC/>A)#8EMZ8AGJM_XKbU/T6_>R;;6ag<(VDH
I_L,S9<Qb7Z[:3Ag2E/.bWT[d0TXCDC;A3DG@ECC#bLI3?J^,<3bUJeC]FL2D)3A
9aMDGR@09(_a&5PIX9,I(049RG_NVMfC,2:BMP4KUa?\T3gJG8W&?[Y^U6gC(VZC
\C\JD,TCH#H/H]\5<9>AJc^QXSRgcbaYZ4]N@M.#P]..C\I0WK=O.?/[)=857^HU
?>L]R;cQ>f/KAM/W2V^VfL)^:J;X@ZGF:I0a&;PLX_D+:PN3bb39M<)L2#O-X)\2
QPNM,CN-\?D6L/>4-,d)[+TD]Y.B2ZH^C7(ZZ;g;P91M=9:)K_d\S57d^?WgW6@8
;bOS6^C8KVcaKc.=\0164d+M^8MV)E>ZYV,VE?0H-V7M>BT</6d[#7@:fFcb\4\Y
bV0&d6S9fH[/SSRdKHD#EN-Qc0PC.C2Wg3?_8L#YXd5\eR#dS0D\(NN[e<IVJ9H?
=M@,?1JYe+V+7QP_?ADKMf1_K-ce0P7Qb31?8/3(M?T8bD)P+H/H7/AM;,CJ=:YS
PNB.(=UM6T2G;d;dEdbS&HG;D[(d5eTV13G=Pg6>L,MZ5M,&C)a7,cD?KF^P2I5W
&RJ0,?c8[7[<:QP(75bF+e]3&d:IU1f2gZJV-:L4Yd81?#,.3#6XB>ES]5MQ2;c-
]QCB9;07C?YD)()6K=V?3W3-15/VMS8()[)H.<9A6bCNW)8]:GA-C,,f8(b<23Ef
U:.XeCP.0E/[ALGS1+&/O:]6LEG,&G(HV^#/?@ALDR2C5&])@4_R]X5NI7YVO,?_
I[TDHgJ>V=PV+bI2-#eaD@>&/+-<1?_LGE07_4)NZDIBT^MSb+gCAW#=O\]X4D?C
?2CZ_+Raa0NRS:NNW[8QFO,W\=N/KS&PG+G;IAd@aIH_-M+FMN@OH^:Y_&F,4ORB
.bgE<3agbF:g.@-V(Y?MVU<dfA9H+W3/W2[^L#faWJA1QX-AdB-36Fb^WF-5-+]P
Q;Y&,3Hf(TRMUZTFFYW:a:E:Q=HV+>2DdT?L5\KMA:);:-,aZW0<KPIWa:>Bg89>
GH5PFHT]G+fCI;WFOCc)9aG53U2/:f<HBJ@J/_(faaJe>L;49/OAVEOP]B:?>L))
>c>\144W-cI54A3JU32)UUO@Z^NI[ePcS,1C_)ERYV6\?2644.G(NN+:+>eCFP8G
L+0OCBB2fW1)L4:d?;I&dYH8)UINDVbWFYaME\LWU/>:/=b&GDAGbA[bX=<5AS1@
^Za11PFJb1B/QgaMaCEVX^1)OLH]VbVKGCZ1/@?RC,^+,J,89@43?H&Q)_7_B]La
]]R+O==HJd/6g=#QN;6UE464>/#>X/_?gS#E@aFCI:(b7d(A,>JT#2TXLO=+ObE>
BfNKWX>QY56LRU)F^QA3WO]d2eEgdOf,&0b]-DR)F9DQ+H(K420<e>?P7I8b_)eN
DPU2JS0J\X?#/:Z[gCf,ZX^D[efIZ(>(LCVa:QIX&9Jd]AWSabaOBf[VPT^e_RUT
bbY8IPb#Td-Q?I5&?I-L=\NQESW2:-/P,P[7(g\\ceFaY5SM0=>EKH@<L/XVVELc
,?f(2/M-[>I=@[RES7R6]J?7&VHe)=e:YW7AZ=dTW)BX_f=6PfDAUaV2FP=Ce(c(
7A>RGbJ3>E)RT_f#://H8)f@,d-3YSJ?2BV-a[TDRb=EWb?bRJdg.O-59A#5^4T=
[8PZ_/dVB2-4a>b=L2AEgRAaY^)YS5NHTWW(1cMRLA#K;JW67;d77<aGaagTV2OU
)=1?Y60H,RY<,+:\c9RXK&5T,#_0QJ3X0HDJ>[\2SKK6cHQ:(\7T:KPFMGb?5_J3
(71;gWDG]gI-_TX@ICb5I\OBG-6)N+PeJgKI?_(g2:20^124a.Rf<8)5/f78QV\G
J_)N-O/e;?8088CabO@B;PTO>.Z30GbM&<Zf?Pe6RL<NX&+8K5FN45/+db3UaT@=
0>=MH4g^deg\.57&K@OQ\S:.F<_VKbU3667_?HK97JP<N4Rce>KOeQ13AB6<E:4?
G,W5;/_;&P1W,5HL1:))+[V@a,E1K/VINNLO]WRW=O/ZDHeeJYN/C<aG/f0590eF
DNaS-S2/;R/.>KbEEH:7MW<&gX,5.A)e5B1<M2]D5O@5(TZCg<ceb&NNC5[+J<;Q
0^Ub3E9fGI-&0VK5;9-1];b^5EG&8JHgBX16X>.(??SQ]H#D&>,J3.KdfBGUSY@e
B=;LU^[._YIT\-&<bEG&ad:MPZO.\-LJGG+&;<,I)U1-5bE[2VdM+02d3bYOH1X+
b5M-Y(e.S),YMSg\A7IK>KGS4IGC<,8+NS49c)8fPS&M]6e9e6/OPV#V8,_HQgd9
1#JBW0X\G9@e6U/L@IDRF12(4S@,2SCc/-=TZb]10V_6&G#M=M9IBI&R_21P;2Ed
7O_S/c\00-M_4F,QI.4?3[XX+FUU6BV(g64A+;_GL5BR?[1dT)UIYADJY6G=?1,X
+dVS\NAU#PG55bH0W1)Mc;<Q(O=J\Mf/JE>U+P/7@[GOD&S^.a:#2JP4@eIT0&CF
+?a2LTb2-@^+L<_J1We@B\eLNEFN>&@C;/eGZ+=3<&7U8gQf2bX9>INT(+6;MM>;
>,/:<;a3&)17+0P:C;A9f9U)UP<R<)A2;#^FN2_L/XY\3MDab]JQ7@d5P:QESf5Q
e7(,b?&L@3X2I69]]D^,JY5b)<Cb.30>J+@+YQ(RC5Q@(A.-I,G)a77W(R5L_R/+
E:3?Qa:5CNLUEg&c=UH8Gf4Zbc8?/ZQ(.)[(YePB=,d<#dHS98O)Ka<8-6N1LC(8
<V?X#]R3ER2<PRWTaT>@H4\b.#MPNe=^:&eA1P98[\;D)5)CDX[T>]>6[,CXZP44
+eO_U+I56)S(DR8C43@&2dCaH?d>Qee=6,bd&7aB>HRP>7DJ?[@\;D8G_fY:Z<F^
;MBM4[L^?-N:ae^4E8:^GI/2\LOcfPYA9Z3.IZ&^F8^MbE(+F,RD:C\Ab)-=V\__
BFYOC(69cYDXI)1V3V2bJ3GfTDZTga^#cU2=a)SbM4VR,Kb/=ES_DBGICgMPc(Ba
O27,dR>bdW1TEQPEcK?3LDa81d(X<<N&DIO0S_B@=HPVOd9R4>-1]+]]U96;\UKc
cPJLe2E,(C/);3MUfVR8HPa#T,&KK0?V#T8ZY9D>UE[6HQ@O7dRRZ;8983E@(39T
/>C5+GfZJbKc:>T93[82=I>JO83bUAJ1JKgLFQB0_KT)RQG0I_@A&KbDeUP:[C\1
+JKA+A0F>d)PfB3[S7JMP^DfD8S[^0LMJ0+I?-@_&c773[)BReZ^:9JZ:fPgYC4[
U0Q+4AFH&2,d.<C2=]/Vc;PC>2cG33F4OE+B-#+dfSKQE.]<@M\G59]^8ML],C;T
+TR<=D8H^-B&X1.[I03I6eS)<aE0MIW@e+e,BgB0L,&T,9NHR7JGGc_HWAI>^g@g
Jc^RH\V7G/03.daH&PPe@<gXc<=.3?8+O5QM]]0B+06S8/T0;6@fR]7E=Fgca_Cc
K.QELN8eE^NNA+X:J.=5WU0\J6FUdSOKa[eD.Mg5K<W6aeGUO?I#BfDf6V(2@Q6G
+ZOOFZ3:@4;YT/25BPdCC]CC2R3]BJWB^FD6/:<.H)02YZaKPZFS/C9SLdQWULL9
fcYP8M/DN&e.cb@&-[ESNBf<-H<;WE0_:LSU_(:>+F-OT(J&>J]d?D/365bS8a[]
-,>\NU=2;A=#_X@MaL5@5W7XITDJbDN]A[_W@gA2RV>g#QUGUeg=VI-;cAaE(g][
X@.d@KbIH0TAQ1@,NOD-??-#JE\KNJ9YK.,-[6K;FBITV2<(B#&L6>:,gNE&2HKd
5>&1Ka6:_W^-dA;)Vd=0AZ)?QAHE(1QXBS?P2g8PCVf=VHS[;QBNZb(]:O&7A8K,
T7RZ@N?P);0e2AfM=U+C9=ID,3;7VP3E)RA\<YY,5SE6L._4^XR2]d.+.L#:TaV,
-/Lef8O[JFO2@,B(S[AUUDP-?4c[@Z,>KQeF[8J[e+dO<]f:L8]b#fH@f,+[YW^?
=a_K+\97B;S?8#4fSD-A(A:;EBVQ/a^DdH9&/K@];<9gadF@K\2[P2H@N$
`endprotected
endmodule